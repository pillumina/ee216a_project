
module Neuron_mul_pixel(
 input clk,
 input GlobalReset,
 input [9:0] Timing_ctr,
 input [9:0] Pix_0, // sfix10_En0
 input [9:0] Pix_1, // sfix10_En0
 input [9:0] Pix_2, // sfix10_En0
 input [9:0] Pix_3, // sfix10_En0
 input [9:0] Pix_4, // sfix10_En0
 input [9:0] Pix_5, // sfix10_En0
 input [9:0] Pix_6, // sfix10_En0
 input [9:0] Pix_7, // sfix10_En0
 input [9:0] Pix_8, // sfix10_En0
 input [9:0] Pix_9, // sfix10_En0
 input [9:0] Pix_10, // sfix10_En0
 input [9:0] Pix_11, // sfix10_En0
 input [9:0] Pix_12, // sfix10_En0
 input [9:0] Pix_13, // sfix10_En0
 input [9:0] Pix_14, // sfix10_En0
 input [9:0] Pix_15, // sfix10_En0
 input [9:0] Pix_16, // sfix10_En0
 input [9:0] Pix_17, // sfix10_En0
 input [9:0] Pix_18, // sfix10_En0
 input [9:0] Pix_19, // sfix10_En0
 input [9:0] Pix_20, // sfix10_En0
 input [9:0] Pix_21, // sfix10_En0
 input [9:0] Pix_22, // sfix10_En0
 input [9:0] Pix_23, // sfix10_En0
 input [9:0] Pix_24, // sfix10_En0
 input [9:0] Pix_25, // sfix10_En0
 input [9:0] Pix_26, // sfix10_En0
 input [9:0] Pix_27, // sfix10_En0
 input [9:0] Pix_28, // sfix10_En0
 input [9:0] Pix_29, // sfix10_En0
 input [9:0] Pix_30, // sfix10_En0
 input [9:0] Pix_31, // sfix10_En0
 input [9:0] Pix_32, // sfix10_En0
 input [9:0] Pix_33, // sfix10_En0
 input [9:0] Pix_34, // sfix10_En0
 input [9:0] Pix_35, // sfix10_En0
 input [9:0] Pix_36, // sfix10_En0
 input [9:0] Pix_37, // sfix10_En0
 input [9:0] Pix_38, // sfix10_En0
 input [9:0] Pix_39, // sfix10_En0
 input [9:0] Pix_40, // sfix10_En0
 input [9:0] Pix_41, // sfix10_En0
 input [9:0] Pix_42, // sfix10_En0
 input [9:0] Pix_43, // sfix10_En0
 input [9:0] Pix_44, // sfix10_En0
 input [9:0] Pix_45, // sfix10_En0
 input [9:0] Pix_46, // sfix10_En0
 input [9:0] Pix_47, // sfix10_En0
 input [9:0] Pix_48, // sfix10_En0
 input [9:0] Pix_49, // sfix10_En0
 input [9:0] Pix_50, // sfix10_En0
 input [9:0] Pix_51, // sfix10_En0
 input [9:0] Pix_52, // sfix10_En0
 input [9:0] Pix_53, // sfix10_En0
 input [9:0] Pix_54, // sfix10_En0
 input [9:0] Pix_55, // sfix10_En0
 input [9:0] Pix_56, // sfix10_En0
 input [9:0] Pix_57, // sfix10_En0
 input [9:0] Pix_58, // sfix10_En0
 input [9:0] Pix_59, // sfix10_En0
 input [9:0] Pix_60, // sfix10_En0
 input [9:0] Pix_61, // sfix10_En0
 input [9:0] Pix_62, // sfix10_En0
 input [9:0] Pix_63, // sfix10_En0
 input [9:0] Pix_64, // sfix10_En0
 input [9:0] Pix_65, // sfix10_En0
 input [9:0] Pix_66, // sfix10_En0
 input [9:0] Pix_67, // sfix10_En0
 input [9:0] Pix_68, // sfix10_En0
 input [9:0] Pix_69, // sfix10_En0
 input [9:0] Pix_70, // sfix10_En0
 input [9:0] Pix_71, // sfix10_En0
 input [9:0] Pix_72, // sfix10_En0
 input [9:0] Pix_73, // sfix10_En0
 input [9:0] Pix_74, // sfix10_En0
 input [9:0] Pix_75, // sfix10_En0
 input [9:0] Pix_76, // sfix10_En0
 input [9:0] Pix_77, // sfix10_En0
 input [9:0] Pix_78, // sfix10_En0
 input [9:0] Pix_79, // sfix10_En0
 input [9:0] Pix_80, // sfix10_En0
 input [9:0] Pix_81, // sfix10_En0
 input [9:0] Pix_82, // sfix10_En0
 input [9:0] Pix_83, // sfix10_En0
 input [9:0] Pix_84, // sfix10_En0
 input [9:0] Pix_85, // sfix10_En0
 input [9:0] Pix_86, // sfix10_En0
 input [9:0] Pix_87, // sfix10_En0
 input [9:0] Pix_88, // sfix10_En0
 input [9:0] Pix_89, // sfix10_En0
 input [9:0] Pix_90, // sfix10_En0
 input [9:0] Pix_91, // sfix10_En0
 input [9:0] Pix_92, // sfix10_En0
 input [9:0] Pix_93, // sfix10_En0
 input [9:0] Pix_94, // sfix10_En0
 input [9:0] Pix_95, // sfix10_En0
 input [9:0] Pix_96, // sfix10_En0
 input [9:0] Pix_97, // sfix10_En0
 input [9:0] Pix_98, // sfix10_En0
 input [9:0] Pix_99, // sfix10_En0
 input [9:0] Pix_100, // sfix10_En0
 input [9:0] Pix_101, // sfix10_En0
 input [9:0] Pix_102, // sfix10_En0
 input [9:0] Pix_103, // sfix10_En0
 input [9:0] Pix_104, // sfix10_En0
 input [9:0] Pix_105, // sfix10_En0
 input [9:0] Pix_106, // sfix10_En0
 input [9:0] Pix_107, // sfix10_En0
 input [9:0] Pix_108, // sfix10_En0
 input [9:0] Pix_109, // sfix10_En0
 input [9:0] Pix_110, // sfix10_En0
 input [9:0] Pix_111, // sfix10_En0
 input [9:0] Pix_112, // sfix10_En0
 input [9:0] Pix_113, // sfix10_En0
 input [9:0] Pix_114, // sfix10_En0
 input [9:0] Pix_115, // sfix10_En0
 input [9:0] Pix_116, // sfix10_En0
 input [9:0] Pix_117, // sfix10_En0
 input [9:0] Pix_118, // sfix10_En0
 input [9:0] Pix_119, // sfix10_En0
 input [9:0] Pix_120, // sfix10_En0
 input [9:0] Pix_121, // sfix10_En0
 input [9:0] Pix_122, // sfix10_En0
 input [9:0] Pix_123, // sfix10_En0
 input [9:0] Pix_124, // sfix10_En0
 input [9:0] Pix_125, // sfix10_En0
 input [9:0] Pix_126, // sfix10_En0
 input [9:0] Pix_127, // sfix10_En0
 input [9:0] Pix_128, // sfix10_En0
 input [9:0] Pix_129, // sfix10_En0
 input [9:0] Pix_130, // sfix10_En0
 input [9:0] Pix_131, // sfix10_En0
 input [9:0] Pix_132, // sfix10_En0
 input [9:0] Pix_133, // sfix10_En0
 input [9:0] Pix_134, // sfix10_En0
 input [9:0] Pix_135, // sfix10_En0
 input [9:0] Pix_136, // sfix10_En0
 input [9:0] Pix_137, // sfix10_En0
 input [9:0] Pix_138, // sfix10_En0
 input [9:0] Pix_139, // sfix10_En0
 input [9:0] Pix_140, // sfix10_En0
 input [9:0] Pix_141, // sfix10_En0
 input [9:0] Pix_142, // sfix10_En0
 input [9:0] Pix_143, // sfix10_En0
 input [9:0] Pix_144, // sfix10_En0
 input [9:0] Pix_145, // sfix10_En0
 input [9:0] Pix_146, // sfix10_En0
 input [9:0] Pix_147, // sfix10_En0
 input [9:0] Pix_148, // sfix10_En0
 input [9:0] Pix_149, // sfix10_En0
 input [9:0] Pix_150, // sfix10_En0
 input [9:0] Pix_151, // sfix10_En0
 input [9:0] Pix_152, // sfix10_En0
 input [9:0] Pix_153, // sfix10_En0
 input [9:0] Pix_154, // sfix10_En0
 input [9:0] Pix_155, // sfix10_En0
 input [9:0] Pix_156, // sfix10_En0
 input [9:0] Pix_157, // sfix10_En0
 input [9:0] Pix_158, // sfix10_En0
 input [9:0] Pix_159, // sfix10_En0
 input [9:0] Pix_160, // sfix10_En0
 input [9:0] Pix_161, // sfix10_En0
 input [9:0] Pix_162, // sfix10_En0
 input [9:0] Pix_163, // sfix10_En0
 input [9:0] Pix_164, // sfix10_En0
 input [9:0] Pix_165, // sfix10_En0
 input [9:0] Pix_166, // sfix10_En0
 input [9:0] Pix_167, // sfix10_En0
 input [9:0] Pix_168, // sfix10_En0
 input [9:0] Pix_169, // sfix10_En0
 input [9:0] Pix_170, // sfix10_En0
 input [9:0] Pix_171, // sfix10_En0
 input [9:0] Pix_172, // sfix10_En0
 input [9:0] Pix_173, // sfix10_En0
 input [9:0] Pix_174, // sfix10_En0
 input [9:0] Pix_175, // sfix10_En0
 input [9:0] Pix_176, // sfix10_En0
 input [9:0] Pix_177, // sfix10_En0
 input [9:0] Pix_178, // sfix10_En0
 input [9:0] Pix_179, // sfix10_En0
 input [9:0] Pix_180, // sfix10_En0
 input [9:0] Pix_181, // sfix10_En0
 input [9:0] Pix_182, // sfix10_En0
 input [9:0] Pix_183, // sfix10_En0
 input [9:0] Pix_184, // sfix10_En0
 input [9:0] Pix_185, // sfix10_En0
 input [9:0] Pix_186, // sfix10_En0
 input [9:0] Pix_187, // sfix10_En0
 input [9:0] Pix_188, // sfix10_En0
 input [9:0] Pix_189, // sfix10_En0
 input [9:0] Pix_190, // sfix10_En0
 input [9:0] Pix_191, // sfix10_En0
 input [9:0] Pix_192, // sfix10_En0
 input [9:0] Pix_193, // sfix10_En0
 input [9:0] Pix_194, // sfix10_En0
 input [9:0] Pix_195, // sfix10_En0
 input [9:0] Pix_196, // sfix10_En0
 input [9:0] Pix_197, // sfix10_En0
 input [9:0] Pix_198, // sfix10_En0
 input [9:0] Pix_199, // sfix10_En0
 input [9:0] Pix_200, // sfix10_En0
 input [9:0] Pix_201, // sfix10_En0
 input [9:0] Pix_202, // sfix10_En0
 input [9:0] Pix_203, // sfix10_En0
 input [9:0] Pix_204, // sfix10_En0
 input [9:0] Pix_205, // sfix10_En0
 input [9:0] Pix_206, // sfix10_En0
 input [9:0] Pix_207, // sfix10_En0
 input [9:0] Pix_208, // sfix10_En0
 input [9:0] Pix_209, // sfix10_En0
 input [9:0] Pix_210, // sfix10_En0
 input [9:0] Pix_211, // sfix10_En0
 input [9:0] Pix_212, // sfix10_En0
 input [9:0] Pix_213, // sfix10_En0
 input [9:0] Pix_214, // sfix10_En0
 input [9:0] Pix_215, // sfix10_En0
 input [9:0] Pix_216, // sfix10_En0
 input [9:0] Pix_217, // sfix10_En0
 input [9:0] Pix_218, // sfix10_En0
 input [9:0] Pix_219, // sfix10_En0
 input [9:0] Pix_220, // sfix10_En0
 input [9:0] Pix_221, // sfix10_En0
 input [9:0] Pix_222, // sfix10_En0
 input [9:0] Pix_223, // sfix10_En0
 input [9:0] Pix_224, // sfix10_En0
 input [9:0] Pix_225, // sfix10_En0
 input [9:0] Pix_226, // sfix10_En0
 input [9:0] Pix_227, // sfix10_En0
 input [9:0] Pix_228, // sfix10_En0
 input [9:0] Pix_229, // sfix10_En0
 input [9:0] Pix_230, // sfix10_En0
 input [9:0] Pix_231, // sfix10_En0
 input [9:0] Pix_232, // sfix10_En0
 input [9:0] Pix_233, // sfix10_En0
 input [9:0] Pix_234, // sfix10_En0
 input [9:0] Pix_235, // sfix10_En0
 input [9:0] Pix_236, // sfix10_En0
 input [9:0] Pix_237, // sfix10_En0
 input [9:0] Pix_238, // sfix10_En0
 input [9:0] Pix_239, // sfix10_En0
 input [9:0] Pix_240, // sfix10_En0
 input [9:0] Pix_241, // sfix10_En0
 input [9:0] Pix_242, // sfix10_En0
 input [9:0] Pix_243, // sfix10_En0
 input [9:0] Pix_244, // sfix10_En0
 input [9:0] Pix_245, // sfix10_En0
 input [9:0] Pix_246, // sfix10_En0
 input [9:0] Pix_247, // sfix10_En0
 input [9:0] Pix_248, // sfix10_En0
 input [9:0] Pix_249, // sfix10_En0
 input [9:0] Pix_250, // sfix10_En0
 input [9:0] Pix_251, // sfix10_En0
 input [9:0] Pix_252, // sfix10_En0
 input [9:0] Pix_253, // sfix10_En0
 input [9:0] Pix_254, // sfix10_En0
 input [9:0] Pix_255, // sfix10_En0
 input [9:0] Pix_256, // sfix10_En0
 input [9:0] Pix_257, // sfix10_En0
 input [9:0] Pix_258, // sfix10_En0
 input [9:0] Pix_259, // sfix10_En0
 input [9:0] Pix_260, // sfix10_En0
 input [9:0] Pix_261, // sfix10_En0
 input [9:0] Pix_262, // sfix10_En0
 input [9:0] Pix_263, // sfix10_En0
 input [9:0] Pix_264, // sfix10_En0
 input [9:0] Pix_265, // sfix10_En0
 input [9:0] Pix_266, // sfix10_En0
 input [9:0] Pix_267, // sfix10_En0
 input [9:0] Pix_268, // sfix10_En0
 input [9:0] Pix_269, // sfix10_En0
 input [9:0] Pix_270, // sfix10_En0
 input [9:0] Pix_271, // sfix10_En0
 input [9:0] Pix_272, // sfix10_En0
 input [9:0] Pix_273, // sfix10_En0
 input [9:0] Pix_274, // sfix10_En0
 input [9:0] Pix_275, // sfix10_En0
 input [9:0] Pix_276, // sfix10_En0
 input [9:0] Pix_277, // sfix10_En0
 input [9:0] Pix_278, // sfix10_En0
 input [9:0] Pix_279, // sfix10_En0
 input [9:0] Pix_280, // sfix10_En0
 input [9:0] Pix_281, // sfix10_En0
 input [9:0] Pix_282, // sfix10_En0
 input [9:0] Pix_283, // sfix10_En0
 input [9:0] Pix_284, // sfix10_En0
 input [9:0] Pix_285, // sfix10_En0
 input [9:0] Pix_286, // sfix10_En0
 input [9:0] Pix_287, // sfix10_En0
 input [9:0] Pix_288, // sfix10_En0
 input [9:0] Pix_289, // sfix10_En0
 input [9:0] Pix_290, // sfix10_En0
 input [9:0] Pix_291, // sfix10_En0
 input [9:0] Pix_292, // sfix10_En0
 input [9:0] Pix_293, // sfix10_En0
 input [9:0] Pix_294, // sfix10_En0
 input [9:0] Pix_295, // sfix10_En0
 input [9:0] Pix_296, // sfix10_En0
 input [9:0] Pix_297, // sfix10_En0
 input [9:0] Pix_298, // sfix10_En0
 input [9:0] Pix_299, // sfix10_En0
 input [9:0] Pix_300, // sfix10_En0
 input [9:0] Pix_301, // sfix10_En0
 input [9:0] Pix_302, // sfix10_En0
 input [9:0] Pix_303, // sfix10_En0
 input [9:0] Pix_304, // sfix10_En0
 input [9:0] Pix_305, // sfix10_En0
 input [9:0] Pix_306, // sfix10_En0
 input [9:0] Pix_307, // sfix10_En0
 input [9:0] Pix_308, // sfix10_En0
 input [9:0] Pix_309, // sfix10_En0
 input [9:0] Pix_310, // sfix10_En0
 input [9:0] Pix_311, // sfix10_En0
 input [9:0] Pix_312, // sfix10_En0
 input [9:0] Pix_313, // sfix10_En0
 input [9:0] Pix_314, // sfix10_En0
 input [9:0] Pix_315, // sfix10_En0
 input [9:0] Pix_316, // sfix10_En0
 input [9:0] Pix_317, // sfix10_En0
 input [9:0] Pix_318, // sfix10_En0
 input [9:0] Pix_319, // sfix10_En0
 input [9:0] Pix_320, // sfix10_En0
 input [9:0] Pix_321, // sfix10_En0
 input [9:0] Pix_322, // sfix10_En0
 input [9:0] Pix_323, // sfix10_En0
 input [9:0] Pix_324, // sfix10_En0
 input [9:0] Pix_325, // sfix10_En0
 input [9:0] Pix_326, // sfix10_En0
 input [9:0] Pix_327, // sfix10_En0
 input [9:0] Pix_328, // sfix10_En0
 input [9:0] Pix_329, // sfix10_En0
 input [9:0] Pix_330, // sfix10_En0
 input [9:0] Pix_331, // sfix10_En0
 input [9:0] Pix_332, // sfix10_En0
 input [9:0] Pix_333, // sfix10_En0
 input [9:0] Pix_334, // sfix10_En0
 input [9:0] Pix_335, // sfix10_En0
 input [9:0] Pix_336, // sfix10_En0
 input [9:0] Pix_337, // sfix10_En0
 input [9:0] Pix_338, // sfix10_En0
 input [9:0] Pix_339, // sfix10_En0
 input [9:0] Pix_340, // sfix10_En0
 input [9:0] Pix_341, // sfix10_En0
 input [9:0] Pix_342, // sfix10_En0
 input [9:0] Pix_343, // sfix10_En0
 input [9:0] Pix_344, // sfix10_En0
 input [9:0] Pix_345, // sfix10_En0
 input [9:0] Pix_346, // sfix10_En0
 input [9:0] Pix_347, // sfix10_En0
 input [9:0] Pix_348, // sfix10_En0
 input [9:0] Pix_349, // sfix10_En0
 input [9:0] Pix_350, // sfix10_En0
 input [9:0] Pix_351, // sfix10_En0
 input [9:0] Pix_352, // sfix10_En0
 input [9:0] Pix_353, // sfix10_En0
 input [9:0] Pix_354, // sfix10_En0
 input [9:0] Pix_355, // sfix10_En0
 input [9:0] Pix_356, // sfix10_En0
 input [9:0] Pix_357, // sfix10_En0
 input [9:0] Pix_358, // sfix10_En0
 input [9:0] Pix_359, // sfix10_En0
 input [9:0] Pix_360, // sfix10_En0
 input [9:0] Pix_361, // sfix10_En0
 input [9:0] Pix_362, // sfix10_En0
 input [9:0] Pix_363, // sfix10_En0
 input [9:0] Pix_364, // sfix10_En0
 input [9:0] Pix_365, // sfix10_En0
 input [9:0] Pix_366, // sfix10_En0
 input [9:0] Pix_367, // sfix10_En0
 input [9:0] Pix_368, // sfix10_En0
 input [9:0] Pix_369, // sfix10_En0
 input [9:0] Pix_370, // sfix10_En0
 input [9:0] Pix_371, // sfix10_En0
 input [9:0] Pix_372, // sfix10_En0
 input [9:0] Pix_373, // sfix10_En0
 input [9:0] Pix_374, // sfix10_En0
 input [9:0] Pix_375, // sfix10_En0
 input [9:0] Pix_376, // sfix10_En0
 input [9:0] Pix_377, // sfix10_En0
 input [9:0] Pix_378, // sfix10_En0
 input [9:0] Pix_379, // sfix10_En0
 input [9:0] Pix_380, // sfix10_En0
 input [9:0] Pix_381, // sfix10_En0
 input [9:0] Pix_382, // sfix10_En0
 input [9:0] Pix_383, // sfix10_En0
 input [9:0] Pix_384, // sfix10_En0
 input [9:0] Pix_385, // sfix10_En0
 input [9:0] Pix_386, // sfix10_En0
 input [9:0] Pix_387, // sfix10_En0
 input [9:0] Pix_388, // sfix10_En0
 input [9:0] Pix_389, // sfix10_En0
 input [9:0] Pix_390, // sfix10_En0
 input [9:0] Pix_391, // sfix10_En0
 input [9:0] Pix_392, // sfix10_En0
 input [9:0] Pix_393, // sfix10_En0
 input [9:0] Pix_394, // sfix10_En0
 input [9:0] Pix_395, // sfix10_En0
 input [9:0] Pix_396, // sfix10_En0
 input [9:0] Pix_397, // sfix10_En0
 input [9:0] Pix_398, // sfix10_En0
 input [9:0] Pix_399, // sfix10_En0
 input [9:0] Pix_400, // sfix10_En0
 input [9:0] Pix_401, // sfix10_En0
 input [9:0] Pix_402, // sfix10_En0
 input [9:0] Pix_403, // sfix10_En0
 input [9:0] Pix_404, // sfix10_En0
 input [9:0] Pix_405, // sfix10_En0
 input [9:0] Pix_406, // sfix10_En0
 input [9:0] Pix_407, // sfix10_En0
 input [9:0] Pix_408, // sfix10_En0
 input [9:0] Pix_409, // sfix10_En0
 input [9:0] Pix_410, // sfix10_En0
 input [9:0] Pix_411, // sfix10_En0
 input [9:0] Pix_412, // sfix10_En0
 input [9:0] Pix_413, // sfix10_En0
 input [9:0] Pix_414, // sfix10_En0
 input [9:0] Pix_415, // sfix10_En0
 input [9:0] Pix_416, // sfix10_En0
 input [9:0] Pix_417, // sfix10_En0
 input [9:0] Pix_418, // sfix10_En0
 input [9:0] Pix_419, // sfix10_En0
 input [9:0] Pix_420, // sfix10_En0
 input [9:0] Pix_421, // sfix10_En0
 input [9:0] Pix_422, // sfix10_En0
 input [9:0] Pix_423, // sfix10_En0
 input [9:0] Pix_424, // sfix10_En0
 input [9:0] Pix_425, // sfix10_En0
 input [9:0] Pix_426, // sfix10_En0
 input [9:0] Pix_427, // sfix10_En0
 input [9:0] Pix_428, // sfix10_En0
 input [9:0] Pix_429, // sfix10_En0
 input [9:0] Pix_430, // sfix10_En0
 input [9:0] Pix_431, // sfix10_En0
 input [9:0] Pix_432, // sfix10_En0
 input [9:0] Pix_433, // sfix10_En0
 input [9:0] Pix_434, // sfix10_En0
 input [9:0] Pix_435, // sfix10_En0
 input [9:0] Pix_436, // sfix10_En0
 input [9:0] Pix_437, // sfix10_En0
 input [9:0] Pix_438, // sfix10_En0
 input [9:0] Pix_439, // sfix10_En0
 input [9:0] Pix_440, // sfix10_En0
 input [9:0] Pix_441, // sfix10_En0
 input [9:0] Pix_442, // sfix10_En0
 input [9:0] Pix_443, // sfix10_En0
 input [9:0] Pix_444, // sfix10_En0
 input [9:0] Pix_445, // sfix10_En0
 input [9:0] Pix_446, // sfix10_En0
 input [9:0] Pix_447, // sfix10_En0
 input [9:0] Pix_448, // sfix10_En0
 input [9:0] Pix_449, // sfix10_En0
 input [9:0] Pix_450, // sfix10_En0
 input [9:0] Pix_451, // sfix10_En0
 input [9:0] Pix_452, // sfix10_En0
 input [9:0] Pix_453, // sfix10_En0
 input [9:0] Pix_454, // sfix10_En0
 input [9:0] Pix_455, // sfix10_En0
 input [9:0] Pix_456, // sfix10_En0
 input [9:0] Pix_457, // sfix10_En0
 input [9:0] Pix_458, // sfix10_En0
 input [9:0] Pix_459, // sfix10_En0
 input [9:0] Pix_460, // sfix10_En0
 input [9:0] Pix_461, // sfix10_En0
 input [9:0] Pix_462, // sfix10_En0
 input [9:0] Pix_463, // sfix10_En0
 input [9:0] Pix_464, // sfix10_En0
 input [9:0] Pix_465, // sfix10_En0
 input [9:0] Pix_466, // sfix10_En0
 input [9:0] Pix_467, // sfix10_En0
 input [9:0] Pix_468, // sfix10_En0
 input [9:0] Pix_469, // sfix10_En0
 input [9:0] Pix_470, // sfix10_En0
 input [9:0] Pix_471, // sfix10_En0
 input [9:0] Pix_472, // sfix10_En0
 input [9:0] Pix_473, // sfix10_En0
 input [9:0] Pix_474, // sfix10_En0
 input [9:0] Pix_475, // sfix10_En0
 input [9:0] Pix_476, // sfix10_En0
 input [9:0] Pix_477, // sfix10_En0
 input [9:0] Pix_478, // sfix10_En0
 input [9:0] Pix_479, // sfix10_En0
 input [9:0] Pix_480, // sfix10_En0
 input [9:0] Pix_481, // sfix10_En0
 input [9:0] Pix_482, // sfix10_En0
 input [9:0] Pix_483, // sfix10_En0
 input [9:0] Pix_484, // sfix10_En0
 input [9:0] Pix_485, // sfix10_En0
 input [9:0] Pix_486, // sfix10_En0
 input [9:0] Pix_487, // sfix10_En0
 input [9:0] Pix_488, // sfix10_En0
 input [9:0] Pix_489, // sfix10_En0
 input [9:0] Pix_490, // sfix10_En0
 input [9:0] Pix_491, // sfix10_En0
 input [9:0] Pix_492, // sfix10_En0
 input [9:0] Pix_493, // sfix10_En0
 input [9:0] Pix_494, // sfix10_En0
 input [9:0] Pix_495, // sfix10_En0
 input [9:0] Pix_496, // sfix10_En0
 input [9:0] Pix_497, // sfix10_En0
 input [9:0] Pix_498, // sfix10_En0
 input [9:0] Pix_499, // sfix10_En0
 input [9:0] Pix_500, // sfix10_En0
 input [9:0] Pix_501, // sfix10_En0
 input [9:0] Pix_502, // sfix10_En0
 input [9:0] Pix_503, // sfix10_En0
 input [9:0] Pix_504, // sfix10_En0
 input [9:0] Pix_505, // sfix10_En0
 input [9:0] Pix_506, // sfix10_En0
 input [9:0] Pix_507, // sfix10_En0
 input [9:0] Pix_508, // sfix10_En0
 input [9:0] Pix_509, // sfix10_En0
 input [9:0] Pix_510, // sfix10_En0
 input [9:0] Pix_511, // sfix10_En0
 input [9:0] Pix_512, // sfix10_En0
 input [9:0] Pix_513, // sfix10_En0
 input [9:0] Pix_514, // sfix10_En0
 input [9:0] Pix_515, // sfix10_En0
 input [9:0] Pix_516, // sfix10_En0
 input [9:0] Pix_517, // sfix10_En0
 input [9:0] Pix_518, // sfix10_En0
 input [9:0] Pix_519, // sfix10_En0
 input [9:0] Pix_520, // sfix10_En0
 input [9:0] Pix_521, // sfix10_En0
 input [9:0] Pix_522, // sfix10_En0
 input [9:0] Pix_523, // sfix10_En0
 input [9:0] Pix_524, // sfix10_En0
 input [9:0] Pix_525, // sfix10_En0
 input [9:0] Pix_526, // sfix10_En0
 input [9:0] Pix_527, // sfix10_En0
 input [9:0] Pix_528, // sfix10_En0
 input [9:0] Pix_529, // sfix10_En0
 input [9:0] Pix_530, // sfix10_En0
 input [9:0] Pix_531, // sfix10_En0
 input [9:0] Pix_532, // sfix10_En0
 input [9:0] Pix_533, // sfix10_En0
 input [9:0] Pix_534, // sfix10_En0
 input [9:0] Pix_535, // sfix10_En0
 input [9:0] Pix_536, // sfix10_En0
 input [9:0] Pix_537, // sfix10_En0
 input [9:0] Pix_538, // sfix10_En0
 input [9:0] Pix_539, // sfix10_En0
 input [9:0] Pix_540, // sfix10_En0
 input [9:0] Pix_541, // sfix10_En0
 input [9:0] Pix_542, // sfix10_En0
 input [9:0] Pix_543, // sfix10_En0
 input [9:0] Pix_544, // sfix10_En0
 input [9:0] Pix_545, // sfix10_En0
 input [9:0] Pix_546, // sfix10_En0
 input [9:0] Pix_547, // sfix10_En0
 input [9:0] Pix_548, // sfix10_En0
 input [9:0] Pix_549, // sfix10_En0
 input [9:0] Pix_550, // sfix10_En0
 input [9:0] Pix_551, // sfix10_En0
 input [9:0] Pix_552, // sfix10_En0
 input [9:0] Pix_553, // sfix10_En0
 input [9:0] Pix_554, // sfix10_En0
 input [9:0] Pix_555, // sfix10_En0
 input [9:0] Pix_556, // sfix10_En0
 input [9:0] Pix_557, // sfix10_En0
 input [9:0] Pix_558, // sfix10_En0
 input [9:0] Pix_559, // sfix10_En0
 input [9:0] Pix_560, // sfix10_En0
 input [9:0] Pix_561, // sfix10_En0
 input [9:0] Pix_562, // sfix10_En0
 input [9:0] Pix_563, // sfix10_En0
 input [9:0] Pix_564, // sfix10_En0
 input [9:0] Pix_565, // sfix10_En0
 input [9:0] Pix_566, // sfix10_En0
 input [9:0] Pix_567, // sfix10_En0
 input [9:0] Pix_568, // sfix10_En0
 input [9:0] Pix_569, // sfix10_En0
 input [9:0] Pix_570, // sfix10_En0
 input [9:0] Pix_571, // sfix10_En0
 input [9:0] Pix_572, // sfix10_En0
 input [9:0] Pix_573, // sfix10_En0
 input [9:0] Pix_574, // sfix10_En0
 input [9:0] Pix_575, // sfix10_En0
 input [9:0] Pix_576, // sfix10_En0
 input [9:0] Pix_577, // sfix10_En0
 input [9:0] Pix_578, // sfix10_En0
 input [9:0] Pix_579, // sfix10_En0
 input [9:0] Pix_580, // sfix10_En0
 input [9:0] Pix_581, // sfix10_En0
 input [9:0] Pix_582, // sfix10_En0
 input [9:0] Pix_583, // sfix10_En0
 input [9:0] Pix_584, // sfix10_En0
 input [9:0] Pix_585, // sfix10_En0
 input [9:0] Pix_586, // sfix10_En0
 input [9:0] Pix_587, // sfix10_En0
 input [9:0] Pix_588, // sfix10_En0
 input [9:0] Pix_589, // sfix10_En0
 input [9:0] Pix_590, // sfix10_En0
 input [9:0] Pix_591, // sfix10_En0
 input [9:0] Pix_592, // sfix10_En0
 input [9:0] Pix_593, // sfix10_En0
 input [9:0] Pix_594, // sfix10_En0
 input [9:0] Pix_595, // sfix10_En0
 input [9:0] Pix_596, // sfix10_En0
 input [9:0] Pix_597, // sfix10_En0
 input [9:0] Pix_598, // sfix10_En0
 input [9:0] Pix_599, // sfix10_En0
 input [9:0] Pix_600, // sfix10_En0
 input [9:0] Pix_601, // sfix10_En0
 input [9:0] Pix_602, // sfix10_En0
 input [9:0] Pix_603, // sfix10_En0
 input [9:0] Pix_604, // sfix10_En0
 input [9:0] Pix_605, // sfix10_En0
 input [9:0] Pix_606, // sfix10_En0
 input [9:0] Pix_607, // sfix10_En0
 input [9:0] Pix_608, // sfix10_En0
 input [9:0] Pix_609, // sfix10_En0
 input [9:0] Pix_610, // sfix10_En0
 input [9:0] Pix_611, // sfix10_En0
 input [9:0] Pix_612, // sfix10_En0
 input [9:0] Pix_613, // sfix10_En0
 input [9:0] Pix_614, // sfix10_En0
 input [9:0] Pix_615, // sfix10_En0
 input [9:0] Pix_616, // sfix10_En0
 input [9:0] Pix_617, // sfix10_En0
 input [9:0] Pix_618, // sfix10_En0
 input [9:0] Pix_619, // sfix10_En0
 input [9:0] Pix_620, // sfix10_En0
 input [9:0] Pix_621, // sfix10_En0
 input [9:0] Pix_622, // sfix10_En0
 input [9:0] Pix_623, // sfix10_En0
 input [9:0] Pix_624, // sfix10_En0
 input [9:0] Pix_625, // sfix10_En0
 input [9:0] Pix_626, // sfix10_En0
 input [9:0] Pix_627, // sfix10_En0
 input [9:0] Pix_628, // sfix10_En0
 input [9:0] Pix_629, // sfix10_En0
 input [9:0] Pix_630, // sfix10_En0
 input [9:0] Pix_631, // sfix10_En0
 input [9:0] Pix_632, // sfix10_En0
 input [9:0] Pix_633, // sfix10_En0
 input [9:0] Pix_634, // sfix10_En0
 input [9:0] Pix_635, // sfix10_En0
 input [9:0] Pix_636, // sfix10_En0
 input [9:0] Pix_637, // sfix10_En0
 input [9:0] Pix_638, // sfix10_En0
 input [9:0] Pix_639, // sfix10_En0
 input [9:0] Pix_640, // sfix10_En0
 input [9:0] Pix_641, // sfix10_En0
 input [9:0] Pix_642, // sfix10_En0
 input [9:0] Pix_643, // sfix10_En0
 input [9:0] Pix_644, // sfix10_En0
 input [9:0] Pix_645, // sfix10_En0
 input [9:0] Pix_646, // sfix10_En0
 input [9:0] Pix_647, // sfix10_En0
 input [9:0] Pix_648, // sfix10_En0
 input [9:0] Pix_649, // sfix10_En0
 input [9:0] Pix_650, // sfix10_En0
 input [9:0] Pix_651, // sfix10_En0
 input [9:0] Pix_652, // sfix10_En0
 input [9:0] Pix_653, // sfix10_En0
 input [9:0] Pix_654, // sfix10_En0
 input [9:0] Pix_655, // sfix10_En0
 input [9:0] Pix_656, // sfix10_En0
 input [9:0] Pix_657, // sfix10_En0
 input [9:0] Pix_658, // sfix10_En0
 input [9:0] Pix_659, // sfix10_En0
 input [9:0] Pix_660, // sfix10_En0
 input [9:0] Pix_661, // sfix10_En0
 input [9:0] Pix_662, // sfix10_En0
 input [9:0] Pix_663, // sfix10_En0
 input [9:0] Pix_664, // sfix10_En0
 input [9:0] Pix_665, // sfix10_En0
 input [9:0] Pix_666, // sfix10_En0
 input [9:0] Pix_667, // sfix10_En0
 input [9:0] Pix_668, // sfix10_En0
 input [9:0] Pix_669, // sfix10_En0
 input [9:0] Pix_670, // sfix10_En0
 input [9:0] Pix_671, // sfix10_En0
 input [9:0] Pix_672, // sfix10_En0
 input [9:0] Pix_673, // sfix10_En0
 input [9:0] Pix_674, // sfix10_En0
 input [9:0] Pix_675, // sfix10_En0
 input [9:0] Pix_676, // sfix10_En0
 input [9:0] Pix_677, // sfix10_En0
 input [9:0] Pix_678, // sfix10_En0
 input [9:0] Pix_679, // sfix10_En0
 input [9:0] Pix_680, // sfix10_En0
 input [9:0] Pix_681, // sfix10_En0
 input [9:0] Pix_682, // sfix10_En0
 input [9:0] Pix_683, // sfix10_En0
 input [9:0] Pix_684, // sfix10_En0
 input [9:0] Pix_685, // sfix10_En0
 input [9:0] Pix_686, // sfix10_En0
 input [9:0] Pix_687, // sfix10_En0
 input [9:0] Pix_688, // sfix10_En0
 input [9:0] Pix_689, // sfix10_En0
 input [9:0] Pix_690, // sfix10_En0
 input [9:0] Pix_691, // sfix10_En0
 input [9:0] Pix_692, // sfix10_En0
 input [9:0] Pix_693, // sfix10_En0
 input [9:0] Pix_694, // sfix10_En0
 input [9:0] Pix_695, // sfix10_En0
 input [9:0] Pix_696, // sfix10_En0
 input [9:0] Pix_697, // sfix10_En0
 input [9:0] Pix_698, // sfix10_En0
 input [9:0] Pix_699, // sfix10_En0
 input [9:0] Pix_700, // sfix10_En0
 input [9:0] Pix_701, // sfix10_En0
 input [9:0] Pix_702, // sfix10_En0
 input [9:0] Pix_703, // sfix10_En0
 input [9:0] Pix_704, // sfix10_En0
 input [9:0] Pix_705, // sfix10_En0
 input [9:0] Pix_706, // sfix10_En0
 input [9:0] Pix_707, // sfix10_En0
 input [9:0] Pix_708, // sfix10_En0
 input [9:0] Pix_709, // sfix10_En0
 input [9:0] Pix_710, // sfix10_En0
 input [9:0] Pix_711, // sfix10_En0
 input [9:0] Pix_712, // sfix10_En0
 input [9:0] Pix_713, // sfix10_En0
 input [9:0] Pix_714, // sfix10_En0
 input [9:0] Pix_715, // sfix10_En0
 input [9:0] Pix_716, // sfix10_En0
 input [9:0] Pix_717, // sfix10_En0
 input [9:0] Pix_718, // sfix10_En0
 input [9:0] Pix_719, // sfix10_En0
 input [9:0] Pix_720, // sfix10_En0
 input [9:0] Pix_721, // sfix10_En0
 input [9:0] Pix_722, // sfix10_En0
 input [9:0] Pix_723, // sfix10_En0
 input [9:0] Pix_724, // sfix10_En0
 input [9:0] Pix_725, // sfix10_En0
 input [9:0] Pix_726, // sfix10_En0
 input [9:0] Pix_727, // sfix10_En0
 input [9:0] Pix_728, // sfix10_En0
 input [9:0] Pix_729, // sfix10_En0
 input [9:0] Pix_730, // sfix10_En0
 input [9:0] Pix_731, // sfix10_En0
 input [9:0] Pix_732, // sfix10_En0
 input [9:0] Pix_733, // sfix10_En0
 input [9:0] Pix_734, // sfix10_En0
 input [9:0] Pix_735, // sfix10_En0
 input [9:0] Pix_736, // sfix10_En0
 input [9:0] Pix_737, // sfix10_En0
 input [9:0] Pix_738, // sfix10_En0
 input [9:0] Pix_739, // sfix10_En0
 input [9:0] Pix_740, // sfix10_En0
 input [9:0] Pix_741, // sfix10_En0
 input [9:0] Pix_742, // sfix10_En0
 input [9:0] Pix_743, // sfix10_En0
 input [9:0] Pix_744, // sfix10_En0
 input [9:0] Pix_745, // sfix10_En0
 input [9:0] Pix_746, // sfix10_En0
 input [9:0] Pix_747, // sfix10_En0
 input [9:0] Pix_748, // sfix10_En0
 input [9:0] Pix_749, // sfix10_En0
 input [9:0] Pix_750, // sfix10_En0
 input [9:0] Pix_751, // sfix10_En0
 input [9:0] Pix_752, // sfix10_En0
 input [9:0] Pix_753, // sfix10_En0
 input [9:0] Pix_754, // sfix10_En0
 input [9:0] Pix_755, // sfix10_En0
 input [9:0] Pix_756, // sfix10_En0
 input [9:0] Pix_757, // sfix10_En0
 input [9:0] Pix_758, // sfix10_En0
 input [9:0] Pix_759, // sfix10_En0
 input [9:0] Pix_760, // sfix10_En0
 input [9:0] Pix_761, // sfix10_En0
 input [9:0] Pix_762, // sfix10_En0
 input [9:0] Pix_763, // sfix10_En0
 input [9:0] Pix_764, // sfix10_En0
 input [9:0] Pix_765, // sfix10_En0
 input [9:0] Pix_766, // sfix10_En0
 input [9:0] Pix_767, // sfix10_En0
 input [9:0] Pix_768, // sfix10_En0
 input [9:0] Pix_769, // sfix10_En0
 input [9:0] Pix_770, // sfix10_En0
 input [9:0] Pix_771, // sfix10_En0
 input [9:0] Pix_772, // sfix10_En0
 input [9:0] Pix_773, // sfix10_En0
 input [9:0] Pix_774, // sfix10_En0
 input [9:0] Pix_775, // sfix10_En0
 input [9:0] Pix_776, // sfix10_En0
 input [9:0] Pix_777, // sfix10_En0
 input [9:0] Pix_778, // sfix10_En0
 input [9:0] Pix_779, // sfix10_En0
 input [9:0] Pix_780, // sfix10_En0
 input [9:0] Pix_781, // sfix10_En0
 input [9:0] Pix_782, // sfix10_En0
 input [9:0] Pix_783, // sfix10_En0
 input [9:0] Pix_784, // sfix10_En0
 output reg [9:0] neuron_0_mul_0_p,
 output reg [9:0] neuron_0_mul_1_p,
 output reg [9:0] neuron_0_mul_2_p,
 output reg [9:0] neuron_0_mul_3_p,
 output reg [9:0] neuron_0_mul_4_p,
 output reg [9:0] neuron_0_mul_5_p,
 output reg [9:0] neuron_0_mul_6_p,
 output reg [9:0] neuron_0_mul_7_p,
 output reg [9:0] neuron_0_mul_8_p,
 output reg [9:0] neuron_0_mul_9_p,
 output reg [9:0] neuron_0_mul_10_p,
 output reg [9:0] neuron_0_mul_11_p,
 output reg [9:0] neuron_0_mul_12_p,
 output reg [9:0] neuron_0_mul_13_p,
 output reg [9:0] neuron_0_mul_14_p,
 output reg [9:0] neuron_0_mul_15_p,
 output reg [9:0] neuron_0_mul_16_p,
 output reg [9:0] neuron_0_mul_17_p,
 output reg [9:0] neuron_0_mul_18_p,
 output reg [9:0] neuron_0_mul_19_p,
 output reg [9:0] neuron_0_mul_20_p,
 output reg [9:0] neuron_0_mul_21_p,
 output reg [9:0] neuron_0_mul_22_p,
 output reg [9:0] neuron_0_mul_23_p,
 output reg [9:0] neuron_0_mul_24_p,
 output reg [9:0] neuron_0_mul_25_p,
 output reg [9:0] neuron_0_mul_26_p,
 output reg [9:0] neuron_0_mul_27_p,
 output reg [9:0] neuron_1_mul_0_p,
 output reg [9:0] neuron_1_mul_1_p,
 output reg [9:0] neuron_1_mul_2_p,
 output reg [9:0] neuron_1_mul_3_p,
 output reg [9:0] neuron_1_mul_4_p,
 output reg [9:0] neuron_1_mul_5_p,
 output reg [9:0] neuron_1_mul_6_p,
 output reg [9:0] neuron_1_mul_7_p,
 output reg [9:0] neuron_1_mul_8_p,
 output reg [9:0] neuron_1_mul_9_p,
 output reg [9:0] neuron_1_mul_10_p,
 output reg [9:0] neuron_1_mul_11_p,
 output reg [9:0] neuron_1_mul_12_p,
 output reg [9:0] neuron_1_mul_13_p,
 output reg [9:0] neuron_1_mul_14_p,
 output reg [9:0] neuron_1_mul_15_p,
 output reg [9:0] neuron_1_mul_16_p,
 output reg [9:0] neuron_1_mul_17_p,
 output reg [9:0] neuron_1_mul_18_p,
 output reg [9:0] neuron_1_mul_19_p,
 output reg [9:0] neuron_1_mul_20_p,
 output reg [9:0] neuron_1_mul_21_p,
 output reg [9:0] neuron_1_mul_22_p,
 output reg [9:0] neuron_1_mul_23_p,
 output reg [9:0] neuron_1_mul_24_p,
 output reg [9:0] neuron_1_mul_25_p,
 output reg [9:0] neuron_1_mul_26_p,
 output reg [9:0] neuron_1_mul_27_p,
 output reg [9:0] neuron_2_mul_0_p,
 output reg [9:0] neuron_2_mul_1_p,
 output reg [9:0] neuron_2_mul_2_p,
 output reg [9:0] neuron_2_mul_3_p,
 output reg [9:0] neuron_2_mul_4_p,
 output reg [9:0] neuron_2_mul_5_p,
 output reg [9:0] neuron_2_mul_6_p,
 output reg [9:0] neuron_2_mul_7_p,
 output reg [9:0] neuron_2_mul_8_p,
 output reg [9:0] neuron_2_mul_9_p,
 output reg [9:0] neuron_2_mul_10_p,
 output reg [9:0] neuron_2_mul_11_p,
 output reg [9:0] neuron_2_mul_12_p,
 output reg [9:0] neuron_2_mul_13_p,
 output reg [9:0] neuron_2_mul_14_p,
 output reg [9:0] neuron_2_mul_15_p,
 output reg [9:0] neuron_2_mul_16_p,
 output reg [9:0] neuron_2_mul_17_p,
 output reg [9:0] neuron_2_mul_18_p,
 output reg [9:0] neuron_2_mul_19_p,
 output reg [9:0] neuron_2_mul_20_p,
 output reg [9:0] neuron_2_mul_21_p,
 output reg [9:0] neuron_2_mul_22_p,
 output reg [9:0] neuron_2_mul_23_p,
 output reg [9:0] neuron_2_mul_24_p,
 output reg [9:0] neuron_2_mul_25_p,
 output reg [9:0] neuron_2_mul_26_p,
 output reg [9:0] neuron_2_mul_27_p,
 output reg [9:0] neuron_3_mul_0_p,
 output reg [9:0] neuron_3_mul_1_p,
 output reg [9:0] neuron_3_mul_2_p,
 output reg [9:0] neuron_3_mul_3_p,
 output reg [9:0] neuron_3_mul_4_p,
 output reg [9:0] neuron_3_mul_5_p,
 output reg [9:0] neuron_3_mul_6_p,
 output reg [9:0] neuron_3_mul_7_p,
 output reg [9:0] neuron_3_mul_8_p,
 output reg [9:0] neuron_3_mul_9_p,
 output reg [9:0] neuron_3_mul_10_p,
 output reg [9:0] neuron_3_mul_11_p,
 output reg [9:0] neuron_3_mul_12_p,
 output reg [9:0] neuron_3_mul_13_p,
 output reg [9:0] neuron_3_mul_14_p,
 output reg [9:0] neuron_3_mul_15_p,
 output reg [9:0] neuron_3_mul_16_p,
 output reg [9:0] neuron_3_mul_17_p,
 output reg [9:0] neuron_3_mul_18_p,
 output reg [9:0] neuron_3_mul_19_p,
 output reg [9:0] neuron_3_mul_20_p,
 output reg [9:0] neuron_3_mul_21_p,
 output reg [9:0] neuron_3_mul_22_p,
 output reg [9:0] neuron_3_mul_23_p,
 output reg [9:0] neuron_3_mul_24_p,
 output reg [9:0] neuron_3_mul_25_p,
 output reg [9:0] neuron_3_mul_26_p,
 output reg [9:0] neuron_3_mul_27_p,
 output reg [9:0] neuron_4_mul_0_p,
 output reg [9:0] neuron_4_mul_1_p,
 output reg [9:0] neuron_4_mul_2_p,
 output reg [9:0] neuron_4_mul_3_p,
 output reg [9:0] neuron_4_mul_4_p,
 output reg [9:0] neuron_4_mul_5_p,
 output reg [9:0] neuron_4_mul_6_p,
 output reg [9:0] neuron_4_mul_7_p,
 output reg [9:0] neuron_4_mul_8_p,
 output reg [9:0] neuron_4_mul_9_p,
 output reg [9:0] neuron_4_mul_10_p,
 output reg [9:0] neuron_4_mul_11_p,
 output reg [9:0] neuron_4_mul_12_p,
 output reg [9:0] neuron_4_mul_13_p,
 output reg [9:0] neuron_4_mul_14_p,
 output reg [9:0] neuron_4_mul_15_p,
 output reg [9:0] neuron_4_mul_16_p,
 output reg [9:0] neuron_4_mul_17_p,
 output reg [9:0] neuron_4_mul_18_p,
 output reg [9:0] neuron_4_mul_19_p,
 output reg [9:0] neuron_4_mul_20_p,
 output reg [9:0] neuron_4_mul_21_p,
 output reg [9:0] neuron_4_mul_22_p,
 output reg [9:0] neuron_4_mul_23_p,
 output reg [9:0] neuron_4_mul_24_p,
 output reg [9:0] neuron_4_mul_25_p,
 output reg [9:0] neuron_4_mul_26_p,
 output reg [9:0] neuron_4_mul_27_p,
 output reg [9:0] neuron_5_mul_0_p,
 output reg [9:0] neuron_5_mul_1_p,
 output reg [9:0] neuron_5_mul_2_p,
 output reg [9:0] neuron_5_mul_3_p,
 output reg [9:0] neuron_5_mul_4_p,
 output reg [9:0] neuron_5_mul_5_p,
 output reg [9:0] neuron_5_mul_6_p,
 output reg [9:0] neuron_5_mul_7_p,
 output reg [9:0] neuron_5_mul_8_p,
 output reg [9:0] neuron_5_mul_9_p,
 output reg [9:0] neuron_5_mul_10_p,
 output reg [9:0] neuron_5_mul_11_p,
 output reg [9:0] neuron_5_mul_12_p,
 output reg [9:0] neuron_5_mul_13_p,
 output reg [9:0] neuron_5_mul_14_p,
 output reg [9:0] neuron_5_mul_15_p,
 output reg [9:0] neuron_5_mul_16_p,
 output reg [9:0] neuron_5_mul_17_p,
 output reg [9:0] neuron_5_mul_18_p,
 output reg [9:0] neuron_5_mul_19_p,
 output reg [9:0] neuron_5_mul_20_p,
 output reg [9:0] neuron_5_mul_21_p,
 output reg [9:0] neuron_5_mul_22_p,
 output reg [9:0] neuron_5_mul_23_p,
 output reg [9:0] neuron_5_mul_24_p,
 output reg [9:0] neuron_5_mul_25_p,
 output reg [9:0] neuron_5_mul_26_p,
 output reg [9:0] neuron_5_mul_27_p,
 output reg [9:0] neuron_6_mul_0_p,
 output reg [9:0] neuron_6_mul_1_p,
 output reg [9:0] neuron_6_mul_2_p,
 output reg [9:0] neuron_6_mul_3_p,
 output reg [9:0] neuron_6_mul_4_p,
 output reg [9:0] neuron_6_mul_5_p,
 output reg [9:0] neuron_6_mul_6_p,
 output reg [9:0] neuron_6_mul_7_p,
 output reg [9:0] neuron_6_mul_8_p,
 output reg [9:0] neuron_6_mul_9_p,
 output reg [9:0] neuron_6_mul_10_p,
 output reg [9:0] neuron_6_mul_11_p,
 output reg [9:0] neuron_6_mul_12_p,
 output reg [9:0] neuron_6_mul_13_p,
 output reg [9:0] neuron_6_mul_14_p,
 output reg [9:0] neuron_6_mul_15_p,
 output reg [9:0] neuron_6_mul_16_p,
 output reg [9:0] neuron_6_mul_17_p,
 output reg [9:0] neuron_6_mul_18_p,
 output reg [9:0] neuron_6_mul_19_p,
 output reg [9:0] neuron_6_mul_20_p,
 output reg [9:0] neuron_6_mul_21_p,
 output reg [9:0] neuron_6_mul_22_p,
 output reg [9:0] neuron_6_mul_23_p,
 output reg [9:0] neuron_6_mul_24_p,
 output reg [9:0] neuron_6_mul_25_p,
 output reg [9:0] neuron_6_mul_26_p,
 output reg [9:0] neuron_6_mul_27_p,
 output reg [9:0] neuron_7_mul_0_p,
 output reg [9:0] neuron_7_mul_1_p,
 output reg [9:0] neuron_7_mul_2_p,
 output reg [9:0] neuron_7_mul_3_p,
 output reg [9:0] neuron_7_mul_4_p,
 output reg [9:0] neuron_7_mul_5_p,
 output reg [9:0] neuron_7_mul_6_p,
 output reg [9:0] neuron_7_mul_7_p,
 output reg [9:0] neuron_7_mul_8_p,
 output reg [9:0] neuron_7_mul_9_p,
 output reg [9:0] neuron_7_mul_10_p,
 output reg [9:0] neuron_7_mul_11_p,
 output reg [9:0] neuron_7_mul_12_p,
 output reg [9:0] neuron_7_mul_13_p,
 output reg [9:0] neuron_7_mul_14_p,
 output reg [9:0] neuron_7_mul_15_p,
 output reg [9:0] neuron_7_mul_16_p,
 output reg [9:0] neuron_7_mul_17_p,
 output reg [9:0] neuron_7_mul_18_p,
 output reg [9:0] neuron_7_mul_19_p,
 output reg [9:0] neuron_7_mul_20_p,
 output reg [9:0] neuron_7_mul_21_p,
 output reg [9:0] neuron_7_mul_22_p,
 output reg [9:0] neuron_7_mul_23_p,
 output reg [9:0] neuron_7_mul_24_p,
 output reg [9:0] neuron_7_mul_25_p,
 output reg [9:0] neuron_7_mul_26_p,
 output reg [9:0] neuron_7_mul_27_p,
 output reg [9:0] neuron_8_mul_0_p,
 output reg [9:0] neuron_8_mul_1_p,
 output reg [9:0] neuron_8_mul_2_p,
 output reg [9:0] neuron_8_mul_3_p,
 output reg [9:0] neuron_8_mul_4_p,
 output reg [9:0] neuron_8_mul_5_p,
 output reg [9:0] neuron_8_mul_6_p,
 output reg [9:0] neuron_8_mul_7_p,
 output reg [9:0] neuron_8_mul_8_p,
 output reg [9:0] neuron_8_mul_9_p,
 output reg [9:0] neuron_8_mul_10_p,
 output reg [9:0] neuron_8_mul_11_p,
 output reg [9:0] neuron_8_mul_12_p,
 output reg [9:0] neuron_8_mul_13_p,
 output reg [9:0] neuron_8_mul_14_p,
 output reg [9:0] neuron_8_mul_15_p,
 output reg [9:0] neuron_8_mul_16_p,
 output reg [9:0] neuron_8_mul_17_p,
 output reg [9:0] neuron_8_mul_18_p,
 output reg [9:0] neuron_8_mul_19_p,
 output reg [9:0] neuron_8_mul_20_p,
 output reg [9:0] neuron_8_mul_21_p,
 output reg [9:0] neuron_8_mul_22_p,
 output reg [9:0] neuron_8_mul_23_p,
 output reg [9:0] neuron_8_mul_24_p,
 output reg [9:0] neuron_8_mul_25_p,
 output reg [9:0] neuron_8_mul_26_p,
 output reg [9:0] neuron_8_mul_27_p,
 output reg [9:0] neuron_9_mul_0_p,
 output reg [9:0] neuron_9_mul_1_p,
 output reg [9:0] neuron_9_mul_2_p,
 output reg [9:0] neuron_9_mul_3_p,
 output reg [9:0] neuron_9_mul_4_p,
 output reg [9:0] neuron_9_mul_5_p,
 output reg [9:0] neuron_9_mul_6_p,
 output reg [9:0] neuron_9_mul_7_p,
 output reg [9:0] neuron_9_mul_8_p,
 output reg [9:0] neuron_9_mul_9_p,
 output reg [9:0] neuron_9_mul_10_p,
 output reg [9:0] neuron_9_mul_11_p,
 output reg [9:0] neuron_9_mul_12_p,
 output reg [9:0] neuron_9_mul_13_p,
 output reg [9:0] neuron_9_mul_14_p,
 output reg [9:0] neuron_9_mul_15_p,
 output reg [9:0] neuron_9_mul_16_p,
 output reg [9:0] neuron_9_mul_17_p,
 output reg [9:0] neuron_9_mul_18_p,
 output reg [9:0] neuron_9_mul_19_p,
 output reg [9:0] neuron_9_mul_20_p,
 output reg [9:0] neuron_9_mul_21_p,
 output reg [9:0] neuron_9_mul_22_p,
 output reg [9:0] neuron_9_mul_23_p,
 output reg [9:0] neuron_9_mul_24_p,
 output reg [9:0] neuron_9_mul_25_p,
 output reg [9:0] neuron_9_mul_26_p,
 output reg [9:0] neuron_9_mul_27_p

);

// For pixels, the blocks below need to be duplicated 27 times
always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_0_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_0_p <= Pix_0;
    10'd1:  neuron_0_mul_0_p <= Pix_1;
    10'd2:  neuron_0_mul_0_p <= Pix_2;
    10'd3:  neuron_0_mul_0_p <= Pix_3;
    10'd4:  neuron_0_mul_0_p <= Pix_4;
    10'd5:  neuron_0_mul_0_p <= Pix_5;
    10'd6:  neuron_0_mul_0_p <= Pix_6;
    10'd7:  neuron_0_mul_0_p <= Pix_7;
    10'd8:  neuron_0_mul_0_p <= Pix_8;
    10'd9:  neuron_0_mul_0_p <= Pix_9;
    10'd10:  neuron_0_mul_0_p <= Pix_10;
    10'd11:  neuron_0_mul_0_p <= Pix_11;
    10'd12:  neuron_0_mul_0_p <= Pix_12;
    10'd13:  neuron_0_mul_0_p <= Pix_13;
    10'd14:  neuron_0_mul_0_p <= Pix_14;
    10'd15:  neuron_0_mul_0_p <= Pix_15;
    10'd16:  neuron_0_mul_0_p <= Pix_16;
    10'd17:  neuron_0_mul_0_p <= Pix_17;
    10'd18:  neuron_0_mul_0_p <= Pix_18;
    10'd19:  neuron_0_mul_0_p <= Pix_19;
    10'd20:  neuron_0_mul_0_p <= Pix_20;
    10'd21:  neuron_0_mul_0_p <= Pix_21;
    10'd22:  neuron_0_mul_0_p <= Pix_22;
    10'd23:  neuron_0_mul_0_p <= Pix_23;
    10'd24:  neuron_0_mul_0_p <= Pix_24;
    10'd25:  neuron_0_mul_0_p <= Pix_25;
    10'd26:  neuron_0_mul_0_p <= Pix_26;
    10'd27:  neuron_0_mul_0_p <= Pix_27;
    default: neuron_0_mul_0_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_1_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_1_p <= Pix_28;
    10'd1:  neuron_0_mul_1_p <= Pix_29;
    10'd2:  neuron_0_mul_1_p <= Pix_30;
    10'd3:  neuron_0_mul_1_p <= Pix_31;
    10'd4:  neuron_0_mul_1_p <= Pix_32;
    10'd5:  neuron_0_mul_1_p <= Pix_33;
    10'd6:  neuron_0_mul_1_p <= Pix_34;
    10'd7:  neuron_0_mul_1_p <= Pix_35;
    10'd8:  neuron_0_mul_1_p <= Pix_36;
    10'd9:  neuron_0_mul_1_p <= Pix_37;
    10'd10:  neuron_0_mul_1_p <= Pix_38;
    10'd11:  neuron_0_mul_1_p <= Pix_39;
    10'd12:  neuron_0_mul_1_p <= Pix_40;
    10'd13:  neuron_0_mul_1_p <= Pix_41;
    10'd14:  neuron_0_mul_1_p <= Pix_42;
    10'd15:  neuron_0_mul_1_p <= Pix_43;
    10'd16:  neuron_0_mul_1_p <= Pix_44;
    10'd17:  neuron_0_mul_1_p <= Pix_45;
    10'd18:  neuron_0_mul_1_p <= Pix_46;
    10'd19:  neuron_0_mul_1_p <= Pix_47;
    10'd20:  neuron_0_mul_1_p <= Pix_48;
    10'd21:  neuron_0_mul_1_p <= Pix_49;
    10'd22:  neuron_0_mul_1_p <= Pix_50;
    10'd23:  neuron_0_mul_1_p <= Pix_51;
    10'd24:  neuron_0_mul_1_p <= Pix_52;
    10'd25:  neuron_0_mul_1_p <= Pix_53;
    10'd26:  neuron_0_mul_1_p <= Pix_54;
    10'd27:  neuron_0_mul_1_p <= Pix_55;
    default: neuron_0_mul_1_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_2_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_2_p <= Pix_56;
    10'd1:  neuron_0_mul_2_p <= Pix_57;
    10'd2:  neuron_0_mul_2_p <= Pix_58;
    10'd3:  neuron_0_mul_2_p <= Pix_59;
    10'd4:  neuron_0_mul_2_p <= Pix_60;
    10'd5:  neuron_0_mul_2_p <= Pix_61;
    10'd6:  neuron_0_mul_2_p <= Pix_62;
    10'd7:  neuron_0_mul_2_p <= Pix_63;
    10'd8:  neuron_0_mul_2_p <= Pix_64;
    10'd9:  neuron_0_mul_2_p <= Pix_65;
    10'd10:  neuron_0_mul_2_p <= Pix_66;
    10'd11:  neuron_0_mul_2_p <= Pix_67;
    10'd12:  neuron_0_mul_2_p <= Pix_68;
    10'd13:  neuron_0_mul_2_p <= Pix_69;
    10'd14:  neuron_0_mul_2_p <= Pix_70;
    10'd15:  neuron_0_mul_2_p <= Pix_71;
    10'd16:  neuron_0_mul_2_p <= Pix_72;
    10'd17:  neuron_0_mul_2_p <= Pix_73;
    10'd18:  neuron_0_mul_2_p <= Pix_74;
    10'd19:  neuron_0_mul_2_p <= Pix_75;
    10'd20:  neuron_0_mul_2_p <= Pix_76;
    10'd21:  neuron_0_mul_2_p <= Pix_77;
    10'd22:  neuron_0_mul_2_p <= Pix_78;
    10'd23:  neuron_0_mul_2_p <= Pix_79;
    10'd24:  neuron_0_mul_2_p <= Pix_80;
    10'd25:  neuron_0_mul_2_p <= Pix_81;
    10'd26:  neuron_0_mul_2_p <= Pix_82;
    10'd27:  neuron_0_mul_2_p <= Pix_83;
    default: neuron_0_mul_2_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_3_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_3_p <= Pix_84;
    10'd1:  neuron_0_mul_3_p <= Pix_85;
    10'd2:  neuron_0_mul_3_p <= Pix_86;
    10'd3:  neuron_0_mul_3_p <= Pix_87;
    10'd4:  neuron_0_mul_3_p <= Pix_88;
    10'd5:  neuron_0_mul_3_p <= Pix_89;
    10'd6:  neuron_0_mul_3_p <= Pix_90;
    10'd7:  neuron_0_mul_3_p <= Pix_91;
    10'd8:  neuron_0_mul_3_p <= Pix_92;
    10'd9:  neuron_0_mul_3_p <= Pix_93;
    10'd10:  neuron_0_mul_3_p <= Pix_94;
    10'd11:  neuron_0_mul_3_p <= Pix_95;
    10'd12:  neuron_0_mul_3_p <= Pix_96;
    10'd13:  neuron_0_mul_3_p <= Pix_97;
    10'd14:  neuron_0_mul_3_p <= Pix_98;
    10'd15:  neuron_0_mul_3_p <= Pix_99;
    10'd16:  neuron_0_mul_3_p <= Pix_100;
    10'd17:  neuron_0_mul_3_p <= Pix_101;
    10'd18:  neuron_0_mul_3_p <= Pix_102;
    10'd19:  neuron_0_mul_3_p <= Pix_103;
    10'd20:  neuron_0_mul_3_p <= Pix_104;
    10'd21:  neuron_0_mul_3_p <= Pix_105;
    10'd22:  neuron_0_mul_3_p <= Pix_106;
    10'd23:  neuron_0_mul_3_p <= Pix_107;
    10'd24:  neuron_0_mul_3_p <= Pix_108;
    10'd25:  neuron_0_mul_3_p <= Pix_109;
    10'd26:  neuron_0_mul_3_p <= Pix_110;
    10'd27:  neuron_0_mul_3_p <= Pix_111;
    default: neuron_0_mul_3_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_4_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_4_p <= Pix_112;
    10'd1:  neuron_0_mul_4_p <= Pix_113;
    10'd2:  neuron_0_mul_4_p <= Pix_114;
    10'd3:  neuron_0_mul_4_p <= Pix_115;
    10'd4:  neuron_0_mul_4_p <= Pix_116;
    10'd5:  neuron_0_mul_4_p <= Pix_117;
    10'd6:  neuron_0_mul_4_p <= Pix_118;
    10'd7:  neuron_0_mul_4_p <= Pix_119;
    10'd8:  neuron_0_mul_4_p <= Pix_120;
    10'd9:  neuron_0_mul_4_p <= Pix_121;
    10'd10:  neuron_0_mul_4_p <= Pix_122;
    10'd11:  neuron_0_mul_4_p <= Pix_123;
    10'd12:  neuron_0_mul_4_p <= Pix_124;
    10'd13:  neuron_0_mul_4_p <= Pix_125;
    10'd14:  neuron_0_mul_4_p <= Pix_126;
    10'd15:  neuron_0_mul_4_p <= Pix_127;
    10'd16:  neuron_0_mul_4_p <= Pix_128;
    10'd17:  neuron_0_mul_4_p <= Pix_129;
    10'd18:  neuron_0_mul_4_p <= Pix_130;
    10'd19:  neuron_0_mul_4_p <= Pix_131;
    10'd20:  neuron_0_mul_4_p <= Pix_132;
    10'd21:  neuron_0_mul_4_p <= Pix_133;
    10'd22:  neuron_0_mul_4_p <= Pix_134;
    10'd23:  neuron_0_mul_4_p <= Pix_135;
    10'd24:  neuron_0_mul_4_p <= Pix_136;
    10'd25:  neuron_0_mul_4_p <= Pix_137;
    10'd26:  neuron_0_mul_4_p <= Pix_138;
    10'd27:  neuron_0_mul_4_p <= Pix_139;
    default: neuron_0_mul_4_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_5_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_5_p <= Pix_140;
    10'd1:  neuron_0_mul_5_p <= Pix_141;
    10'd2:  neuron_0_mul_5_p <= Pix_142;
    10'd3:  neuron_0_mul_5_p <= Pix_143;
    10'd4:  neuron_0_mul_5_p <= Pix_144;
    10'd5:  neuron_0_mul_5_p <= Pix_145;
    10'd6:  neuron_0_mul_5_p <= Pix_146;
    10'd7:  neuron_0_mul_5_p <= Pix_147;
    10'd8:  neuron_0_mul_5_p <= Pix_148;
    10'd9:  neuron_0_mul_5_p <= Pix_149;
    10'd10:  neuron_0_mul_5_p <= Pix_150;
    10'd11:  neuron_0_mul_5_p <= Pix_151;
    10'd12:  neuron_0_mul_5_p <= Pix_152;
    10'd13:  neuron_0_mul_5_p <= Pix_153;
    10'd14:  neuron_0_mul_5_p <= Pix_154;
    10'd15:  neuron_0_mul_5_p <= Pix_155;
    10'd16:  neuron_0_mul_5_p <= Pix_156;
    10'd17:  neuron_0_mul_5_p <= Pix_157;
    10'd18:  neuron_0_mul_5_p <= Pix_158;
    10'd19:  neuron_0_mul_5_p <= Pix_159;
    10'd20:  neuron_0_mul_5_p <= Pix_160;
    10'd21:  neuron_0_mul_5_p <= Pix_161;
    10'd22:  neuron_0_mul_5_p <= Pix_162;
    10'd23:  neuron_0_mul_5_p <= Pix_163;
    10'd24:  neuron_0_mul_5_p <= Pix_164;
    10'd25:  neuron_0_mul_5_p <= Pix_165;
    10'd26:  neuron_0_mul_5_p <= Pix_166;
    10'd27:  neuron_0_mul_5_p <= Pix_167;
    default: neuron_0_mul_5_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_6_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_6_p <= Pix_168;
    10'd1:  neuron_0_mul_6_p <= Pix_169;
    10'd2:  neuron_0_mul_6_p <= Pix_170;
    10'd3:  neuron_0_mul_6_p <= Pix_171;
    10'd4:  neuron_0_mul_6_p <= Pix_172;
    10'd5:  neuron_0_mul_6_p <= Pix_173;
    10'd6:  neuron_0_mul_6_p <= Pix_174;
    10'd7:  neuron_0_mul_6_p <= Pix_175;
    10'd8:  neuron_0_mul_6_p <= Pix_176;
    10'd9:  neuron_0_mul_6_p <= Pix_177;
    10'd10:  neuron_0_mul_6_p <= Pix_178;
    10'd11:  neuron_0_mul_6_p <= Pix_179;
    10'd12:  neuron_0_mul_6_p <= Pix_180;
    10'd13:  neuron_0_mul_6_p <= Pix_181;
    10'd14:  neuron_0_mul_6_p <= Pix_182;
    10'd15:  neuron_0_mul_6_p <= Pix_183;
    10'd16:  neuron_0_mul_6_p <= Pix_184;
    10'd17:  neuron_0_mul_6_p <= Pix_185;
    10'd18:  neuron_0_mul_6_p <= Pix_186;
    10'd19:  neuron_0_mul_6_p <= Pix_187;
    10'd20:  neuron_0_mul_6_p <= Pix_188;
    10'd21:  neuron_0_mul_6_p <= Pix_189;
    10'd22:  neuron_0_mul_6_p <= Pix_190;
    10'd23:  neuron_0_mul_6_p <= Pix_191;
    10'd24:  neuron_0_mul_6_p <= Pix_192;
    10'd25:  neuron_0_mul_6_p <= Pix_193;
    10'd26:  neuron_0_mul_6_p <= Pix_194;
    10'd27:  neuron_0_mul_6_p <= Pix_195;
    default: neuron_0_mul_6_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_7_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_7_p <= Pix_196;
    10'd1:  neuron_0_mul_7_p <= Pix_197;
    10'd2:  neuron_0_mul_7_p <= Pix_198;
    10'd3:  neuron_0_mul_7_p <= Pix_199;
    10'd4:  neuron_0_mul_7_p <= Pix_200;
    10'd5:  neuron_0_mul_7_p <= Pix_201;
    10'd6:  neuron_0_mul_7_p <= Pix_202;
    10'd7:  neuron_0_mul_7_p <= Pix_203;
    10'd8:  neuron_0_mul_7_p <= Pix_204;
    10'd9:  neuron_0_mul_7_p <= Pix_205;
    10'd10:  neuron_0_mul_7_p <= Pix_206;
    10'd11:  neuron_0_mul_7_p <= Pix_207;
    10'd12:  neuron_0_mul_7_p <= Pix_208;
    10'd13:  neuron_0_mul_7_p <= Pix_209;
    10'd14:  neuron_0_mul_7_p <= Pix_210;
    10'd15:  neuron_0_mul_7_p <= Pix_211;
    10'd16:  neuron_0_mul_7_p <= Pix_212;
    10'd17:  neuron_0_mul_7_p <= Pix_213;
    10'd18:  neuron_0_mul_7_p <= Pix_214;
    10'd19:  neuron_0_mul_7_p <= Pix_215;
    10'd20:  neuron_0_mul_7_p <= Pix_216;
    10'd21:  neuron_0_mul_7_p <= Pix_217;
    10'd22:  neuron_0_mul_7_p <= Pix_218;
    10'd23:  neuron_0_mul_7_p <= Pix_219;
    10'd24:  neuron_0_mul_7_p <= Pix_220;
    10'd25:  neuron_0_mul_7_p <= Pix_221;
    10'd26:  neuron_0_mul_7_p <= Pix_222;
    10'd27:  neuron_0_mul_7_p <= Pix_223;
    default: neuron_0_mul_7_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_8_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_8_p <= Pix_224;
    10'd1:  neuron_0_mul_8_p <= Pix_225;
    10'd2:  neuron_0_mul_8_p <= Pix_226;
    10'd3:  neuron_0_mul_8_p <= Pix_227;
    10'd4:  neuron_0_mul_8_p <= Pix_228;
    10'd5:  neuron_0_mul_8_p <= Pix_229;
    10'd6:  neuron_0_mul_8_p <= Pix_230;
    10'd7:  neuron_0_mul_8_p <= Pix_231;
    10'd8:  neuron_0_mul_8_p <= Pix_232;
    10'd9:  neuron_0_mul_8_p <= Pix_233;
    10'd10:  neuron_0_mul_8_p <= Pix_234;
    10'd11:  neuron_0_mul_8_p <= Pix_235;
    10'd12:  neuron_0_mul_8_p <= Pix_236;
    10'd13:  neuron_0_mul_8_p <= Pix_237;
    10'd14:  neuron_0_mul_8_p <= Pix_238;
    10'd15:  neuron_0_mul_8_p <= Pix_239;
    10'd16:  neuron_0_mul_8_p <= Pix_240;
    10'd17:  neuron_0_mul_8_p <= Pix_241;
    10'd18:  neuron_0_mul_8_p <= Pix_242;
    10'd19:  neuron_0_mul_8_p <= Pix_243;
    10'd20:  neuron_0_mul_8_p <= Pix_244;
    10'd21:  neuron_0_mul_8_p <= Pix_245;
    10'd22:  neuron_0_mul_8_p <= Pix_246;
    10'd23:  neuron_0_mul_8_p <= Pix_247;
    10'd24:  neuron_0_mul_8_p <= Pix_248;
    10'd25:  neuron_0_mul_8_p <= Pix_249;
    10'd26:  neuron_0_mul_8_p <= Pix_250;
    10'd27:  neuron_0_mul_8_p <= Pix_251;
    default: neuron_0_mul_8_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_9_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_9_p <= Pix_252;
    10'd1:  neuron_0_mul_9_p <= Pix_253;
    10'd2:  neuron_0_mul_9_p <= Pix_254;
    10'd3:  neuron_0_mul_9_p <= Pix_255;
    10'd4:  neuron_0_mul_9_p <= Pix_256;
    10'd5:  neuron_0_mul_9_p <= Pix_257;
    10'd6:  neuron_0_mul_9_p <= Pix_258;
    10'd7:  neuron_0_mul_9_p <= Pix_259;
    10'd8:  neuron_0_mul_9_p <= Pix_260;
    10'd9:  neuron_0_mul_9_p <= Pix_261;
    10'd10:  neuron_0_mul_9_p <= Pix_262;
    10'd11:  neuron_0_mul_9_p <= Pix_263;
    10'd12:  neuron_0_mul_9_p <= Pix_264;
    10'd13:  neuron_0_mul_9_p <= Pix_265;
    10'd14:  neuron_0_mul_9_p <= Pix_266;
    10'd15:  neuron_0_mul_9_p <= Pix_267;
    10'd16:  neuron_0_mul_9_p <= Pix_268;
    10'd17:  neuron_0_mul_9_p <= Pix_269;
    10'd18:  neuron_0_mul_9_p <= Pix_270;
    10'd19:  neuron_0_mul_9_p <= Pix_271;
    10'd20:  neuron_0_mul_9_p <= Pix_272;
    10'd21:  neuron_0_mul_9_p <= Pix_273;
    10'd22:  neuron_0_mul_9_p <= Pix_274;
    10'd23:  neuron_0_mul_9_p <= Pix_275;
    10'd24:  neuron_0_mul_9_p <= Pix_276;
    10'd25:  neuron_0_mul_9_p <= Pix_277;
    10'd26:  neuron_0_mul_9_p <= Pix_278;
    10'd27:  neuron_0_mul_9_p <= Pix_279;
    default: neuron_0_mul_9_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_10_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_10_p <= Pix_280;
    10'd1:  neuron_0_mul_10_p <= Pix_281;
    10'd2:  neuron_0_mul_10_p <= Pix_282;
    10'd3:  neuron_0_mul_10_p <= Pix_283;
    10'd4:  neuron_0_mul_10_p <= Pix_284;
    10'd5:  neuron_0_mul_10_p <= Pix_285;
    10'd6:  neuron_0_mul_10_p <= Pix_286;
    10'd7:  neuron_0_mul_10_p <= Pix_287;
    10'd8:  neuron_0_mul_10_p <= Pix_288;
    10'd9:  neuron_0_mul_10_p <= Pix_289;
    10'd10:  neuron_0_mul_10_p <= Pix_290;
    10'd11:  neuron_0_mul_10_p <= Pix_291;
    10'd12:  neuron_0_mul_10_p <= Pix_292;
    10'd13:  neuron_0_mul_10_p <= Pix_293;
    10'd14:  neuron_0_mul_10_p <= Pix_294;
    10'd15:  neuron_0_mul_10_p <= Pix_295;
    10'd16:  neuron_0_mul_10_p <= Pix_296;
    10'd17:  neuron_0_mul_10_p <= Pix_297;
    10'd18:  neuron_0_mul_10_p <= Pix_298;
    10'd19:  neuron_0_mul_10_p <= Pix_299;
    10'd20:  neuron_0_mul_10_p <= Pix_300;
    10'd21:  neuron_0_mul_10_p <= Pix_301;
    10'd22:  neuron_0_mul_10_p <= Pix_302;
    10'd23:  neuron_0_mul_10_p <= Pix_303;
    10'd24:  neuron_0_mul_10_p <= Pix_304;
    10'd25:  neuron_0_mul_10_p <= Pix_305;
    10'd26:  neuron_0_mul_10_p <= Pix_306;
    10'd27:  neuron_0_mul_10_p <= Pix_307;
    default: neuron_0_mul_10_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_11_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_11_p <= Pix_308;
    10'd1:  neuron_0_mul_11_p <= Pix_309;
    10'd2:  neuron_0_mul_11_p <= Pix_310;
    10'd3:  neuron_0_mul_11_p <= Pix_311;
    10'd4:  neuron_0_mul_11_p <= Pix_312;
    10'd5:  neuron_0_mul_11_p <= Pix_313;
    10'd6:  neuron_0_mul_11_p <= Pix_314;
    10'd7:  neuron_0_mul_11_p <= Pix_315;
    10'd8:  neuron_0_mul_11_p <= Pix_316;
    10'd9:  neuron_0_mul_11_p <= Pix_317;
    10'd10:  neuron_0_mul_11_p <= Pix_318;
    10'd11:  neuron_0_mul_11_p <= Pix_319;
    10'd12:  neuron_0_mul_11_p <= Pix_320;
    10'd13:  neuron_0_mul_11_p <= Pix_321;
    10'd14:  neuron_0_mul_11_p <= Pix_322;
    10'd15:  neuron_0_mul_11_p <= Pix_323;
    10'd16:  neuron_0_mul_11_p <= Pix_324;
    10'd17:  neuron_0_mul_11_p <= Pix_325;
    10'd18:  neuron_0_mul_11_p <= Pix_326;
    10'd19:  neuron_0_mul_11_p <= Pix_327;
    10'd20:  neuron_0_mul_11_p <= Pix_328;
    10'd21:  neuron_0_mul_11_p <= Pix_329;
    10'd22:  neuron_0_mul_11_p <= Pix_330;
    10'd23:  neuron_0_mul_11_p <= Pix_331;
    10'd24:  neuron_0_mul_11_p <= Pix_332;
    10'd25:  neuron_0_mul_11_p <= Pix_333;
    10'd26:  neuron_0_mul_11_p <= Pix_334;
    10'd27:  neuron_0_mul_11_p <= Pix_335;
    default: neuron_0_mul_11_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_12_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_12_p <= Pix_336;
    10'd1:  neuron_0_mul_12_p <= Pix_337;
    10'd2:  neuron_0_mul_12_p <= Pix_338;
    10'd3:  neuron_0_mul_12_p <= Pix_339;
    10'd4:  neuron_0_mul_12_p <= Pix_340;
    10'd5:  neuron_0_mul_12_p <= Pix_341;
    10'd6:  neuron_0_mul_12_p <= Pix_342;
    10'd7:  neuron_0_mul_12_p <= Pix_343;
    10'd8:  neuron_0_mul_12_p <= Pix_344;
    10'd9:  neuron_0_mul_12_p <= Pix_345;
    10'd10:  neuron_0_mul_12_p <= Pix_346;
    10'd11:  neuron_0_mul_12_p <= Pix_347;
    10'd12:  neuron_0_mul_12_p <= Pix_348;
    10'd13:  neuron_0_mul_12_p <= Pix_349;
    10'd14:  neuron_0_mul_12_p <= Pix_350;
    10'd15:  neuron_0_mul_12_p <= Pix_351;
    10'd16:  neuron_0_mul_12_p <= Pix_352;
    10'd17:  neuron_0_mul_12_p <= Pix_353;
    10'd18:  neuron_0_mul_12_p <= Pix_354;
    10'd19:  neuron_0_mul_12_p <= Pix_355;
    10'd20:  neuron_0_mul_12_p <= Pix_356;
    10'd21:  neuron_0_mul_12_p <= Pix_357;
    10'd22:  neuron_0_mul_12_p <= Pix_358;
    10'd23:  neuron_0_mul_12_p <= Pix_359;
    10'd24:  neuron_0_mul_12_p <= Pix_360;
    10'd25:  neuron_0_mul_12_p <= Pix_361;
    10'd26:  neuron_0_mul_12_p <= Pix_362;
    10'd27:  neuron_0_mul_12_p <= Pix_363;
    default: neuron_0_mul_12_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_13_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_13_p <= Pix_364;
    10'd1:  neuron_0_mul_13_p <= Pix_365;
    10'd2:  neuron_0_mul_13_p <= Pix_366;
    10'd3:  neuron_0_mul_13_p <= Pix_367;
    10'd4:  neuron_0_mul_13_p <= Pix_368;
    10'd5:  neuron_0_mul_13_p <= Pix_369;
    10'd6:  neuron_0_mul_13_p <= Pix_370;
    10'd7:  neuron_0_mul_13_p <= Pix_371;
    10'd8:  neuron_0_mul_13_p <= Pix_372;
    10'd9:  neuron_0_mul_13_p <= Pix_373;
    10'd10:  neuron_0_mul_13_p <= Pix_374;
    10'd11:  neuron_0_mul_13_p <= Pix_375;
    10'd12:  neuron_0_mul_13_p <= Pix_376;
    10'd13:  neuron_0_mul_13_p <= Pix_377;
    10'd14:  neuron_0_mul_13_p <= Pix_378;
    10'd15:  neuron_0_mul_13_p <= Pix_379;
    10'd16:  neuron_0_mul_13_p <= Pix_380;
    10'd17:  neuron_0_mul_13_p <= Pix_381;
    10'd18:  neuron_0_mul_13_p <= Pix_382;
    10'd19:  neuron_0_mul_13_p <= Pix_383;
    10'd20:  neuron_0_mul_13_p <= Pix_384;
    10'd21:  neuron_0_mul_13_p <= Pix_385;
    10'd22:  neuron_0_mul_13_p <= Pix_386;
    10'd23:  neuron_0_mul_13_p <= Pix_387;
    10'd24:  neuron_0_mul_13_p <= Pix_388;
    10'd25:  neuron_0_mul_13_p <= Pix_389;
    10'd26:  neuron_0_mul_13_p <= Pix_390;
    10'd27:  neuron_0_mul_13_p <= Pix_391;
    default: neuron_0_mul_13_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_14_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_14_p <= Pix_392;
    10'd1:  neuron_0_mul_14_p <= Pix_393;
    10'd2:  neuron_0_mul_14_p <= Pix_394;
    10'd3:  neuron_0_mul_14_p <= Pix_395;
    10'd4:  neuron_0_mul_14_p <= Pix_396;
    10'd5:  neuron_0_mul_14_p <= Pix_397;
    10'd6:  neuron_0_mul_14_p <= Pix_398;
    10'd7:  neuron_0_mul_14_p <= Pix_399;
    10'd8:  neuron_0_mul_14_p <= Pix_400;
    10'd9:  neuron_0_mul_14_p <= Pix_401;
    10'd10:  neuron_0_mul_14_p <= Pix_402;
    10'd11:  neuron_0_mul_14_p <= Pix_403;
    10'd12:  neuron_0_mul_14_p <= Pix_404;
    10'd13:  neuron_0_mul_14_p <= Pix_405;
    10'd14:  neuron_0_mul_14_p <= Pix_406;
    10'd15:  neuron_0_mul_14_p <= Pix_407;
    10'd16:  neuron_0_mul_14_p <= Pix_408;
    10'd17:  neuron_0_mul_14_p <= Pix_409;
    10'd18:  neuron_0_mul_14_p <= Pix_410;
    10'd19:  neuron_0_mul_14_p <= Pix_411;
    10'd20:  neuron_0_mul_14_p <= Pix_412;
    10'd21:  neuron_0_mul_14_p <= Pix_413;
    10'd22:  neuron_0_mul_14_p <= Pix_414;
    10'd23:  neuron_0_mul_14_p <= Pix_415;
    10'd24:  neuron_0_mul_14_p <= Pix_416;
    10'd25:  neuron_0_mul_14_p <= Pix_417;
    10'd26:  neuron_0_mul_14_p <= Pix_418;
    10'd27:  neuron_0_mul_14_p <= Pix_419;
    default: neuron_0_mul_14_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_15_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_15_p <= Pix_420;
    10'd1:  neuron_0_mul_15_p <= Pix_421;
    10'd2:  neuron_0_mul_15_p <= Pix_422;
    10'd3:  neuron_0_mul_15_p <= Pix_423;
    10'd4:  neuron_0_mul_15_p <= Pix_424;
    10'd5:  neuron_0_mul_15_p <= Pix_425;
    10'd6:  neuron_0_mul_15_p <= Pix_426;
    10'd7:  neuron_0_mul_15_p <= Pix_427;
    10'd8:  neuron_0_mul_15_p <= Pix_428;
    10'd9:  neuron_0_mul_15_p <= Pix_429;
    10'd10:  neuron_0_mul_15_p <= Pix_430;
    10'd11:  neuron_0_mul_15_p <= Pix_431;
    10'd12:  neuron_0_mul_15_p <= Pix_432;
    10'd13:  neuron_0_mul_15_p <= Pix_433;
    10'd14:  neuron_0_mul_15_p <= Pix_434;
    10'd15:  neuron_0_mul_15_p <= Pix_435;
    10'd16:  neuron_0_mul_15_p <= Pix_436;
    10'd17:  neuron_0_mul_15_p <= Pix_437;
    10'd18:  neuron_0_mul_15_p <= Pix_438;
    10'd19:  neuron_0_mul_15_p <= Pix_439;
    10'd20:  neuron_0_mul_15_p <= Pix_440;
    10'd21:  neuron_0_mul_15_p <= Pix_441;
    10'd22:  neuron_0_mul_15_p <= Pix_442;
    10'd23:  neuron_0_mul_15_p <= Pix_443;
    10'd24:  neuron_0_mul_15_p <= Pix_444;
    10'd25:  neuron_0_mul_15_p <= Pix_445;
    10'd26:  neuron_0_mul_15_p <= Pix_446;
    10'd27:  neuron_0_mul_15_p <= Pix_447;
    default: neuron_0_mul_15_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_16_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_16_p <= Pix_448;
    10'd1:  neuron_0_mul_16_p <= Pix_449;
    10'd2:  neuron_0_mul_16_p <= Pix_450;
    10'd3:  neuron_0_mul_16_p <= Pix_451;
    10'd4:  neuron_0_mul_16_p <= Pix_452;
    10'd5:  neuron_0_mul_16_p <= Pix_453;
    10'd6:  neuron_0_mul_16_p <= Pix_454;
    10'd7:  neuron_0_mul_16_p <= Pix_455;
    10'd8:  neuron_0_mul_16_p <= Pix_456;
    10'd9:  neuron_0_mul_16_p <= Pix_457;
    10'd10:  neuron_0_mul_16_p <= Pix_458;
    10'd11:  neuron_0_mul_16_p <= Pix_459;
    10'd12:  neuron_0_mul_16_p <= Pix_460;
    10'd13:  neuron_0_mul_16_p <= Pix_461;
    10'd14:  neuron_0_mul_16_p <= Pix_462;
    10'd15:  neuron_0_mul_16_p <= Pix_463;
    10'd16:  neuron_0_mul_16_p <= Pix_464;
    10'd17:  neuron_0_mul_16_p <= Pix_465;
    10'd18:  neuron_0_mul_16_p <= Pix_466;
    10'd19:  neuron_0_mul_16_p <= Pix_467;
    10'd20:  neuron_0_mul_16_p <= Pix_468;
    10'd21:  neuron_0_mul_16_p <= Pix_469;
    10'd22:  neuron_0_mul_16_p <= Pix_470;
    10'd23:  neuron_0_mul_16_p <= Pix_471;
    10'd24:  neuron_0_mul_16_p <= Pix_472;
    10'd25:  neuron_0_mul_16_p <= Pix_473;
    10'd26:  neuron_0_mul_16_p <= Pix_474;
    10'd27:  neuron_0_mul_16_p <= Pix_475;
    default: neuron_0_mul_16_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_17_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_17_p <= Pix_476;
    10'd1:  neuron_0_mul_17_p <= Pix_477;
    10'd2:  neuron_0_mul_17_p <= Pix_478;
    10'd3:  neuron_0_mul_17_p <= Pix_479;
    10'd4:  neuron_0_mul_17_p <= Pix_480;
    10'd5:  neuron_0_mul_17_p <= Pix_481;
    10'd6:  neuron_0_mul_17_p <= Pix_482;
    10'd7:  neuron_0_mul_17_p <= Pix_483;
    10'd8:  neuron_0_mul_17_p <= Pix_484;
    10'd9:  neuron_0_mul_17_p <= Pix_485;
    10'd10:  neuron_0_mul_17_p <= Pix_486;
    10'd11:  neuron_0_mul_17_p <= Pix_487;
    10'd12:  neuron_0_mul_17_p <= Pix_488;
    10'd13:  neuron_0_mul_17_p <= Pix_489;
    10'd14:  neuron_0_mul_17_p <= Pix_490;
    10'd15:  neuron_0_mul_17_p <= Pix_491;
    10'd16:  neuron_0_mul_17_p <= Pix_492;
    10'd17:  neuron_0_mul_17_p <= Pix_493;
    10'd18:  neuron_0_mul_17_p <= Pix_494;
    10'd19:  neuron_0_mul_17_p <= Pix_495;
    10'd20:  neuron_0_mul_17_p <= Pix_496;
    10'd21:  neuron_0_mul_17_p <= Pix_497;
    10'd22:  neuron_0_mul_17_p <= Pix_498;
    10'd23:  neuron_0_mul_17_p <= Pix_499;
    10'd24:  neuron_0_mul_17_p <= Pix_500;
    10'd25:  neuron_0_mul_17_p <= Pix_501;
    10'd26:  neuron_0_mul_17_p <= Pix_502;
    10'd27:  neuron_0_mul_17_p <= Pix_503;
    default: neuron_0_mul_17_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_18_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_18_p <= Pix_504;
    10'd1:  neuron_0_mul_18_p <= Pix_505;
    10'd2:  neuron_0_mul_18_p <= Pix_506;
    10'd3:  neuron_0_mul_18_p <= Pix_507;
    10'd4:  neuron_0_mul_18_p <= Pix_508;
    10'd5:  neuron_0_mul_18_p <= Pix_509;
    10'd6:  neuron_0_mul_18_p <= Pix_510;
    10'd7:  neuron_0_mul_18_p <= Pix_511;
    10'd8:  neuron_0_mul_18_p <= Pix_512;
    10'd9:  neuron_0_mul_18_p <= Pix_513;
    10'd10:  neuron_0_mul_18_p <= Pix_514;
    10'd11:  neuron_0_mul_18_p <= Pix_515;
    10'd12:  neuron_0_mul_18_p <= Pix_516;
    10'd13:  neuron_0_mul_18_p <= Pix_517;
    10'd14:  neuron_0_mul_18_p <= Pix_518;
    10'd15:  neuron_0_mul_18_p <= Pix_519;
    10'd16:  neuron_0_mul_18_p <= Pix_520;
    10'd17:  neuron_0_mul_18_p <= Pix_521;
    10'd18:  neuron_0_mul_18_p <= Pix_522;
    10'd19:  neuron_0_mul_18_p <= Pix_523;
    10'd20:  neuron_0_mul_18_p <= Pix_524;
    10'd21:  neuron_0_mul_18_p <= Pix_525;
    10'd22:  neuron_0_mul_18_p <= Pix_526;
    10'd23:  neuron_0_mul_18_p <= Pix_527;
    10'd24:  neuron_0_mul_18_p <= Pix_528;
    10'd25:  neuron_0_mul_18_p <= Pix_529;
    10'd26:  neuron_0_mul_18_p <= Pix_530;
    10'd27:  neuron_0_mul_18_p <= Pix_531;
    default: neuron_0_mul_18_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_19_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_19_p <= Pix_532;
    10'd1:  neuron_0_mul_19_p <= Pix_533;
    10'd2:  neuron_0_mul_19_p <= Pix_534;
    10'd3:  neuron_0_mul_19_p <= Pix_535;
    10'd4:  neuron_0_mul_19_p <= Pix_536;
    10'd5:  neuron_0_mul_19_p <= Pix_537;
    10'd6:  neuron_0_mul_19_p <= Pix_538;
    10'd7:  neuron_0_mul_19_p <= Pix_539;
    10'd8:  neuron_0_mul_19_p <= Pix_540;
    10'd9:  neuron_0_mul_19_p <= Pix_541;
    10'd10:  neuron_0_mul_19_p <= Pix_542;
    10'd11:  neuron_0_mul_19_p <= Pix_543;
    10'd12:  neuron_0_mul_19_p <= Pix_544;
    10'd13:  neuron_0_mul_19_p <= Pix_545;
    10'd14:  neuron_0_mul_19_p <= Pix_546;
    10'd15:  neuron_0_mul_19_p <= Pix_547;
    10'd16:  neuron_0_mul_19_p <= Pix_548;
    10'd17:  neuron_0_mul_19_p <= Pix_549;
    10'd18:  neuron_0_mul_19_p <= Pix_550;
    10'd19:  neuron_0_mul_19_p <= Pix_551;
    10'd20:  neuron_0_mul_19_p <= Pix_552;
    10'd21:  neuron_0_mul_19_p <= Pix_553;
    10'd22:  neuron_0_mul_19_p <= Pix_554;
    10'd23:  neuron_0_mul_19_p <= Pix_555;
    10'd24:  neuron_0_mul_19_p <= Pix_556;
    10'd25:  neuron_0_mul_19_p <= Pix_557;
    10'd26:  neuron_0_mul_19_p <= Pix_558;
    10'd27:  neuron_0_mul_19_p <= Pix_559;
    default: neuron_0_mul_19_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_20_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_20_p <= Pix_560;
    10'd1:  neuron_0_mul_20_p <= Pix_561;
    10'd2:  neuron_0_mul_20_p <= Pix_562;
    10'd3:  neuron_0_mul_20_p <= Pix_563;
    10'd4:  neuron_0_mul_20_p <= Pix_564;
    10'd5:  neuron_0_mul_20_p <= Pix_565;
    10'd6:  neuron_0_mul_20_p <= Pix_566;
    10'd7:  neuron_0_mul_20_p <= Pix_567;
    10'd8:  neuron_0_mul_20_p <= Pix_568;
    10'd9:  neuron_0_mul_20_p <= Pix_569;
    10'd10:  neuron_0_mul_20_p <= Pix_570;
    10'd11:  neuron_0_mul_20_p <= Pix_571;
    10'd12:  neuron_0_mul_20_p <= Pix_572;
    10'd13:  neuron_0_mul_20_p <= Pix_573;
    10'd14:  neuron_0_mul_20_p <= Pix_574;
    10'd15:  neuron_0_mul_20_p <= Pix_575;
    10'd16:  neuron_0_mul_20_p <= Pix_576;
    10'd17:  neuron_0_mul_20_p <= Pix_577;
    10'd18:  neuron_0_mul_20_p <= Pix_578;
    10'd19:  neuron_0_mul_20_p <= Pix_579;
    10'd20:  neuron_0_mul_20_p <= Pix_580;
    10'd21:  neuron_0_mul_20_p <= Pix_581;
    10'd22:  neuron_0_mul_20_p <= Pix_582;
    10'd23:  neuron_0_mul_20_p <= Pix_583;
    10'd24:  neuron_0_mul_20_p <= Pix_584;
    10'd25:  neuron_0_mul_20_p <= Pix_585;
    10'd26:  neuron_0_mul_20_p <= Pix_586;
    10'd27:  neuron_0_mul_20_p <= Pix_587;
    default: neuron_0_mul_20_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_21_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_21_p <= Pix_588;
    10'd1:  neuron_0_mul_21_p <= Pix_589;
    10'd2:  neuron_0_mul_21_p <= Pix_590;
    10'd3:  neuron_0_mul_21_p <= Pix_591;
    10'd4:  neuron_0_mul_21_p <= Pix_592;
    10'd5:  neuron_0_mul_21_p <= Pix_593;
    10'd6:  neuron_0_mul_21_p <= Pix_594;
    10'd7:  neuron_0_mul_21_p <= Pix_595;
    10'd8:  neuron_0_mul_21_p <= Pix_596;
    10'd9:  neuron_0_mul_21_p <= Pix_597;
    10'd10:  neuron_0_mul_21_p <= Pix_598;
    10'd11:  neuron_0_mul_21_p <= Pix_599;
    10'd12:  neuron_0_mul_21_p <= Pix_600;
    10'd13:  neuron_0_mul_21_p <= Pix_601;
    10'd14:  neuron_0_mul_21_p <= Pix_602;
    10'd15:  neuron_0_mul_21_p <= Pix_603;
    10'd16:  neuron_0_mul_21_p <= Pix_604;
    10'd17:  neuron_0_mul_21_p <= Pix_605;
    10'd18:  neuron_0_mul_21_p <= Pix_606;
    10'd19:  neuron_0_mul_21_p <= Pix_607;
    10'd20:  neuron_0_mul_21_p <= Pix_608;
    10'd21:  neuron_0_mul_21_p <= Pix_609;
    10'd22:  neuron_0_mul_21_p <= Pix_610;
    10'd23:  neuron_0_mul_21_p <= Pix_611;
    10'd24:  neuron_0_mul_21_p <= Pix_612;
    10'd25:  neuron_0_mul_21_p <= Pix_613;
    10'd26:  neuron_0_mul_21_p <= Pix_614;
    10'd27:  neuron_0_mul_21_p <= Pix_615;
    default: neuron_0_mul_21_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_22_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_22_p <= Pix_616;
    10'd1:  neuron_0_mul_22_p <= Pix_617;
    10'd2:  neuron_0_mul_22_p <= Pix_618;
    10'd3:  neuron_0_mul_22_p <= Pix_619;
    10'd4:  neuron_0_mul_22_p <= Pix_620;
    10'd5:  neuron_0_mul_22_p <= Pix_621;
    10'd6:  neuron_0_mul_22_p <= Pix_622;
    10'd7:  neuron_0_mul_22_p <= Pix_623;
    10'd8:  neuron_0_mul_22_p <= Pix_624;
    10'd9:  neuron_0_mul_22_p <= Pix_625;
    10'd10:  neuron_0_mul_22_p <= Pix_626;
    10'd11:  neuron_0_mul_22_p <= Pix_627;
    10'd12:  neuron_0_mul_22_p <= Pix_628;
    10'd13:  neuron_0_mul_22_p <= Pix_629;
    10'd14:  neuron_0_mul_22_p <= Pix_630;
    10'd15:  neuron_0_mul_22_p <= Pix_631;
    10'd16:  neuron_0_mul_22_p <= Pix_632;
    10'd17:  neuron_0_mul_22_p <= Pix_633;
    10'd18:  neuron_0_mul_22_p <= Pix_634;
    10'd19:  neuron_0_mul_22_p <= Pix_635;
    10'd20:  neuron_0_mul_22_p <= Pix_636;
    10'd21:  neuron_0_mul_22_p <= Pix_637;
    10'd22:  neuron_0_mul_22_p <= Pix_638;
    10'd23:  neuron_0_mul_22_p <= Pix_639;
    10'd24:  neuron_0_mul_22_p <= Pix_640;
    10'd25:  neuron_0_mul_22_p <= Pix_641;
    10'd26:  neuron_0_mul_22_p <= Pix_642;
    10'd27:  neuron_0_mul_22_p <= Pix_643;
    default: neuron_0_mul_22_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_23_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_23_p <= Pix_644;
    10'd1:  neuron_0_mul_23_p <= Pix_645;
    10'd2:  neuron_0_mul_23_p <= Pix_646;
    10'd3:  neuron_0_mul_23_p <= Pix_647;
    10'd4:  neuron_0_mul_23_p <= Pix_648;
    10'd5:  neuron_0_mul_23_p <= Pix_649;
    10'd6:  neuron_0_mul_23_p <= Pix_650;
    10'd7:  neuron_0_mul_23_p <= Pix_651;
    10'd8:  neuron_0_mul_23_p <= Pix_652;
    10'd9:  neuron_0_mul_23_p <= Pix_653;
    10'd10:  neuron_0_mul_23_p <= Pix_654;
    10'd11:  neuron_0_mul_23_p <= Pix_655;
    10'd12:  neuron_0_mul_23_p <= Pix_656;
    10'd13:  neuron_0_mul_23_p <= Pix_657;
    10'd14:  neuron_0_mul_23_p <= Pix_658;
    10'd15:  neuron_0_mul_23_p <= Pix_659;
    10'd16:  neuron_0_mul_23_p <= Pix_660;
    10'd17:  neuron_0_mul_23_p <= Pix_661;
    10'd18:  neuron_0_mul_23_p <= Pix_662;
    10'd19:  neuron_0_mul_23_p <= Pix_663;
    10'd20:  neuron_0_mul_23_p <= Pix_664;
    10'd21:  neuron_0_mul_23_p <= Pix_665;
    10'd22:  neuron_0_mul_23_p <= Pix_666;
    10'd23:  neuron_0_mul_23_p <= Pix_667;
    10'd24:  neuron_0_mul_23_p <= Pix_668;
    10'd25:  neuron_0_mul_23_p <= Pix_669;
    10'd26:  neuron_0_mul_23_p <= Pix_670;
    10'd27:  neuron_0_mul_23_p <= Pix_671;
    default: neuron_0_mul_23_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_24_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_24_p <= Pix_672;
    10'd1:  neuron_0_mul_24_p <= Pix_673;
    10'd2:  neuron_0_mul_24_p <= Pix_674;
    10'd3:  neuron_0_mul_24_p <= Pix_675;
    10'd4:  neuron_0_mul_24_p <= Pix_676;
    10'd5:  neuron_0_mul_24_p <= Pix_677;
    10'd6:  neuron_0_mul_24_p <= Pix_678;
    10'd7:  neuron_0_mul_24_p <= Pix_679;
    10'd8:  neuron_0_mul_24_p <= Pix_680;
    10'd9:  neuron_0_mul_24_p <= Pix_681;
    10'd10:  neuron_0_mul_24_p <= Pix_682;
    10'd11:  neuron_0_mul_24_p <= Pix_683;
    10'd12:  neuron_0_mul_24_p <= Pix_684;
    10'd13:  neuron_0_mul_24_p <= Pix_685;
    10'd14:  neuron_0_mul_24_p <= Pix_686;
    10'd15:  neuron_0_mul_24_p <= Pix_687;
    10'd16:  neuron_0_mul_24_p <= Pix_688;
    10'd17:  neuron_0_mul_24_p <= Pix_689;
    10'd18:  neuron_0_mul_24_p <= Pix_690;
    10'd19:  neuron_0_mul_24_p <= Pix_691;
    10'd20:  neuron_0_mul_24_p <= Pix_692;
    10'd21:  neuron_0_mul_24_p <= Pix_693;
    10'd22:  neuron_0_mul_24_p <= Pix_694;
    10'd23:  neuron_0_mul_24_p <= Pix_695;
    10'd24:  neuron_0_mul_24_p <= Pix_696;
    10'd25:  neuron_0_mul_24_p <= Pix_697;
    10'd26:  neuron_0_mul_24_p <= Pix_698;
    10'd27:  neuron_0_mul_24_p <= Pix_699;
    default: neuron_0_mul_24_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_25_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_25_p <= Pix_700;
    10'd1:  neuron_0_mul_25_p <= Pix_701;
    10'd2:  neuron_0_mul_25_p <= Pix_702;
    10'd3:  neuron_0_mul_25_p <= Pix_703;
    10'd4:  neuron_0_mul_25_p <= Pix_704;
    10'd5:  neuron_0_mul_25_p <= Pix_705;
    10'd6:  neuron_0_mul_25_p <= Pix_706;
    10'd7:  neuron_0_mul_25_p <= Pix_707;
    10'd8:  neuron_0_mul_25_p <= Pix_708;
    10'd9:  neuron_0_mul_25_p <= Pix_709;
    10'd10:  neuron_0_mul_25_p <= Pix_710;
    10'd11:  neuron_0_mul_25_p <= Pix_711;
    10'd12:  neuron_0_mul_25_p <= Pix_712;
    10'd13:  neuron_0_mul_25_p <= Pix_713;
    10'd14:  neuron_0_mul_25_p <= Pix_714;
    10'd15:  neuron_0_mul_25_p <= Pix_715;
    10'd16:  neuron_0_mul_25_p <= Pix_716;
    10'd17:  neuron_0_mul_25_p <= Pix_717;
    10'd18:  neuron_0_mul_25_p <= Pix_718;
    10'd19:  neuron_0_mul_25_p <= Pix_719;
    10'd20:  neuron_0_mul_25_p <= Pix_720;
    10'd21:  neuron_0_mul_25_p <= Pix_721;
    10'd22:  neuron_0_mul_25_p <= Pix_722;
    10'd23:  neuron_0_mul_25_p <= Pix_723;
    10'd24:  neuron_0_mul_25_p <= Pix_724;
    10'd25:  neuron_0_mul_25_p <= Pix_725;
    10'd26:  neuron_0_mul_25_p <= Pix_726;
    10'd27:  neuron_0_mul_25_p <= Pix_727;
    default: neuron_0_mul_25_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_26_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_26_p <= Pix_728;
    10'd1:  neuron_0_mul_26_p <= Pix_729;
    10'd2:  neuron_0_mul_26_p <= Pix_730;
    10'd3:  neuron_0_mul_26_p <= Pix_731;
    10'd4:  neuron_0_mul_26_p <= Pix_732;
    10'd5:  neuron_0_mul_26_p <= Pix_733;
    10'd6:  neuron_0_mul_26_p <= Pix_734;
    10'd7:  neuron_0_mul_26_p <= Pix_735;
    10'd8:  neuron_0_mul_26_p <= Pix_736;
    10'd9:  neuron_0_mul_26_p <= Pix_737;
    10'd10:  neuron_0_mul_26_p <= Pix_738;
    10'd11:  neuron_0_mul_26_p <= Pix_739;
    10'd12:  neuron_0_mul_26_p <= Pix_740;
    10'd13:  neuron_0_mul_26_p <= Pix_741;
    10'd14:  neuron_0_mul_26_p <= Pix_742;
    10'd15:  neuron_0_mul_26_p <= Pix_743;
    10'd16:  neuron_0_mul_26_p <= Pix_744;
    10'd17:  neuron_0_mul_26_p <= Pix_745;
    10'd18:  neuron_0_mul_26_p <= Pix_746;
    10'd19:  neuron_0_mul_26_p <= Pix_747;
    10'd20:  neuron_0_mul_26_p <= Pix_748;
    10'd21:  neuron_0_mul_26_p <= Pix_749;
    10'd22:  neuron_0_mul_26_p <= Pix_750;
    10'd23:  neuron_0_mul_26_p <= Pix_751;
    10'd24:  neuron_0_mul_26_p <= Pix_752;
    10'd25:  neuron_0_mul_26_p <= Pix_753;
    10'd26:  neuron_0_mul_26_p <= Pix_754;
    10'd27:  neuron_0_mul_26_p <= Pix_755;
    default: neuron_0_mul_26_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_0_mul_27_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_0_mul_27_p <= Pix_756;
    10'd1:  neuron_0_mul_27_p <= Pix_757;
    10'd2:  neuron_0_mul_27_p <= Pix_758;
    10'd3:  neuron_0_mul_27_p <= Pix_759;
    10'd4:  neuron_0_mul_27_p <= Pix_760;
    10'd5:  neuron_0_mul_27_p <= Pix_761;
    10'd6:  neuron_0_mul_27_p <= Pix_762;
    10'd7:  neuron_0_mul_27_p <= Pix_763;
    10'd8:  neuron_0_mul_27_p <= Pix_764;
    10'd9:  neuron_0_mul_27_p <= Pix_765;
    10'd10:  neuron_0_mul_27_p <= Pix_766;
    10'd11:  neuron_0_mul_27_p <= Pix_767;
    10'd12:  neuron_0_mul_27_p <= Pix_768;
    10'd13:  neuron_0_mul_27_p <= Pix_769;
    10'd14:  neuron_0_mul_27_p <= Pix_770;
    10'd15:  neuron_0_mul_27_p <= Pix_771;
    10'd16:  neuron_0_mul_27_p <= Pix_772;
    10'd17:  neuron_0_mul_27_p <= Pix_773;
    10'd18:  neuron_0_mul_27_p <= Pix_774;
    10'd19:  neuron_0_mul_27_p <= Pix_775;
    10'd20:  neuron_0_mul_27_p <= Pix_776;
    10'd21:  neuron_0_mul_27_p <= Pix_777;
    10'd22:  neuron_0_mul_27_p <= Pix_778;
    10'd23:  neuron_0_mul_27_p <= Pix_779;
    10'd24:  neuron_0_mul_27_p <= Pix_780;
    10'd25:  neuron_0_mul_27_p <= Pix_781;
    10'd26:  neuron_0_mul_27_p <= Pix_782;
    10'd27:  neuron_0_mul_27_p <= Pix_783;
    default: neuron_0_mul_27_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_0_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_0_p <= Pix_0;
    10'd1:  neuron_1_mul_0_p <= Pix_1;
    10'd2:  neuron_1_mul_0_p <= Pix_2;
    10'd3:  neuron_1_mul_0_p <= Pix_3;
    10'd4:  neuron_1_mul_0_p <= Pix_4;
    10'd5:  neuron_1_mul_0_p <= Pix_5;
    10'd6:  neuron_1_mul_0_p <= Pix_6;
    10'd7:  neuron_1_mul_0_p <= Pix_7;
    10'd8:  neuron_1_mul_0_p <= Pix_8;
    10'd9:  neuron_1_mul_0_p <= Pix_9;
    10'd10:  neuron_1_mul_0_p <= Pix_10;
    10'd11:  neuron_1_mul_0_p <= Pix_11;
    10'd12:  neuron_1_mul_0_p <= Pix_12;
    10'd13:  neuron_1_mul_0_p <= Pix_13;
    10'd14:  neuron_1_mul_0_p <= Pix_14;
    10'd15:  neuron_1_mul_0_p <= Pix_15;
    10'd16:  neuron_1_mul_0_p <= Pix_16;
    10'd17:  neuron_1_mul_0_p <= Pix_17;
    10'd18:  neuron_1_mul_0_p <= Pix_18;
    10'd19:  neuron_1_mul_0_p <= Pix_19;
    10'd20:  neuron_1_mul_0_p <= Pix_20;
    10'd21:  neuron_1_mul_0_p <= Pix_21;
    10'd22:  neuron_1_mul_0_p <= Pix_22;
    10'd23:  neuron_1_mul_0_p <= Pix_23;
    10'd24:  neuron_1_mul_0_p <= Pix_24;
    10'd25:  neuron_1_mul_0_p <= Pix_25;
    10'd26:  neuron_1_mul_0_p <= Pix_26;
    10'd27:  neuron_1_mul_0_p <= Pix_27;
    default: neuron_1_mul_0_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_1_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_1_p <= Pix_28;
    10'd1:  neuron_1_mul_1_p <= Pix_29;
    10'd2:  neuron_1_mul_1_p <= Pix_30;
    10'd3:  neuron_1_mul_1_p <= Pix_31;
    10'd4:  neuron_1_mul_1_p <= Pix_32;
    10'd5:  neuron_1_mul_1_p <= Pix_33;
    10'd6:  neuron_1_mul_1_p <= Pix_34;
    10'd7:  neuron_1_mul_1_p <= Pix_35;
    10'd8:  neuron_1_mul_1_p <= Pix_36;
    10'd9:  neuron_1_mul_1_p <= Pix_37;
    10'd10:  neuron_1_mul_1_p <= Pix_38;
    10'd11:  neuron_1_mul_1_p <= Pix_39;
    10'd12:  neuron_1_mul_1_p <= Pix_40;
    10'd13:  neuron_1_mul_1_p <= Pix_41;
    10'd14:  neuron_1_mul_1_p <= Pix_42;
    10'd15:  neuron_1_mul_1_p <= Pix_43;
    10'd16:  neuron_1_mul_1_p <= Pix_44;
    10'd17:  neuron_1_mul_1_p <= Pix_45;
    10'd18:  neuron_1_mul_1_p <= Pix_46;
    10'd19:  neuron_1_mul_1_p <= Pix_47;
    10'd20:  neuron_1_mul_1_p <= Pix_48;
    10'd21:  neuron_1_mul_1_p <= Pix_49;
    10'd22:  neuron_1_mul_1_p <= Pix_50;
    10'd23:  neuron_1_mul_1_p <= Pix_51;
    10'd24:  neuron_1_mul_1_p <= Pix_52;
    10'd25:  neuron_1_mul_1_p <= Pix_53;
    10'd26:  neuron_1_mul_1_p <= Pix_54;
    10'd27:  neuron_1_mul_1_p <= Pix_55;
    default: neuron_1_mul_1_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_2_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_2_p <= Pix_56;
    10'd1:  neuron_1_mul_2_p <= Pix_57;
    10'd2:  neuron_1_mul_2_p <= Pix_58;
    10'd3:  neuron_1_mul_2_p <= Pix_59;
    10'd4:  neuron_1_mul_2_p <= Pix_60;
    10'd5:  neuron_1_mul_2_p <= Pix_61;
    10'd6:  neuron_1_mul_2_p <= Pix_62;
    10'd7:  neuron_1_mul_2_p <= Pix_63;
    10'd8:  neuron_1_mul_2_p <= Pix_64;
    10'd9:  neuron_1_mul_2_p <= Pix_65;
    10'd10:  neuron_1_mul_2_p <= Pix_66;
    10'd11:  neuron_1_mul_2_p <= Pix_67;
    10'd12:  neuron_1_mul_2_p <= Pix_68;
    10'd13:  neuron_1_mul_2_p <= Pix_69;
    10'd14:  neuron_1_mul_2_p <= Pix_70;
    10'd15:  neuron_1_mul_2_p <= Pix_71;
    10'd16:  neuron_1_mul_2_p <= Pix_72;
    10'd17:  neuron_1_mul_2_p <= Pix_73;
    10'd18:  neuron_1_mul_2_p <= Pix_74;
    10'd19:  neuron_1_mul_2_p <= Pix_75;
    10'd20:  neuron_1_mul_2_p <= Pix_76;
    10'd21:  neuron_1_mul_2_p <= Pix_77;
    10'd22:  neuron_1_mul_2_p <= Pix_78;
    10'd23:  neuron_1_mul_2_p <= Pix_79;
    10'd24:  neuron_1_mul_2_p <= Pix_80;
    10'd25:  neuron_1_mul_2_p <= Pix_81;
    10'd26:  neuron_1_mul_2_p <= Pix_82;
    10'd27:  neuron_1_mul_2_p <= Pix_83;
    default: neuron_1_mul_2_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_3_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_3_p <= Pix_84;
    10'd1:  neuron_1_mul_3_p <= Pix_85;
    10'd2:  neuron_1_mul_3_p <= Pix_86;
    10'd3:  neuron_1_mul_3_p <= Pix_87;
    10'd4:  neuron_1_mul_3_p <= Pix_88;
    10'd5:  neuron_1_mul_3_p <= Pix_89;
    10'd6:  neuron_1_mul_3_p <= Pix_90;
    10'd7:  neuron_1_mul_3_p <= Pix_91;
    10'd8:  neuron_1_mul_3_p <= Pix_92;
    10'd9:  neuron_1_mul_3_p <= Pix_93;
    10'd10:  neuron_1_mul_3_p <= Pix_94;
    10'd11:  neuron_1_mul_3_p <= Pix_95;
    10'd12:  neuron_1_mul_3_p <= Pix_96;
    10'd13:  neuron_1_mul_3_p <= Pix_97;
    10'd14:  neuron_1_mul_3_p <= Pix_98;
    10'd15:  neuron_1_mul_3_p <= Pix_99;
    10'd16:  neuron_1_mul_3_p <= Pix_100;
    10'd17:  neuron_1_mul_3_p <= Pix_101;
    10'd18:  neuron_1_mul_3_p <= Pix_102;
    10'd19:  neuron_1_mul_3_p <= Pix_103;
    10'd20:  neuron_1_mul_3_p <= Pix_104;
    10'd21:  neuron_1_mul_3_p <= Pix_105;
    10'd22:  neuron_1_mul_3_p <= Pix_106;
    10'd23:  neuron_1_mul_3_p <= Pix_107;
    10'd24:  neuron_1_mul_3_p <= Pix_108;
    10'd25:  neuron_1_mul_3_p <= Pix_109;
    10'd26:  neuron_1_mul_3_p <= Pix_110;
    10'd27:  neuron_1_mul_3_p <= Pix_111;
    default: neuron_1_mul_3_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_4_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_4_p <= Pix_112;
    10'd1:  neuron_1_mul_4_p <= Pix_113;
    10'd2:  neuron_1_mul_4_p <= Pix_114;
    10'd3:  neuron_1_mul_4_p <= Pix_115;
    10'd4:  neuron_1_mul_4_p <= Pix_116;
    10'd5:  neuron_1_mul_4_p <= Pix_117;
    10'd6:  neuron_1_mul_4_p <= Pix_118;
    10'd7:  neuron_1_mul_4_p <= Pix_119;
    10'd8:  neuron_1_mul_4_p <= Pix_120;
    10'd9:  neuron_1_mul_4_p <= Pix_121;
    10'd10:  neuron_1_mul_4_p <= Pix_122;
    10'd11:  neuron_1_mul_4_p <= Pix_123;
    10'd12:  neuron_1_mul_4_p <= Pix_124;
    10'd13:  neuron_1_mul_4_p <= Pix_125;
    10'd14:  neuron_1_mul_4_p <= Pix_126;
    10'd15:  neuron_1_mul_4_p <= Pix_127;
    10'd16:  neuron_1_mul_4_p <= Pix_128;
    10'd17:  neuron_1_mul_4_p <= Pix_129;
    10'd18:  neuron_1_mul_4_p <= Pix_130;
    10'd19:  neuron_1_mul_4_p <= Pix_131;
    10'd20:  neuron_1_mul_4_p <= Pix_132;
    10'd21:  neuron_1_mul_4_p <= Pix_133;
    10'd22:  neuron_1_mul_4_p <= Pix_134;
    10'd23:  neuron_1_mul_4_p <= Pix_135;
    10'd24:  neuron_1_mul_4_p <= Pix_136;
    10'd25:  neuron_1_mul_4_p <= Pix_137;
    10'd26:  neuron_1_mul_4_p <= Pix_138;
    10'd27:  neuron_1_mul_4_p <= Pix_139;
    default: neuron_1_mul_4_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_5_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_5_p <= Pix_140;
    10'd1:  neuron_1_mul_5_p <= Pix_141;
    10'd2:  neuron_1_mul_5_p <= Pix_142;
    10'd3:  neuron_1_mul_5_p <= Pix_143;
    10'd4:  neuron_1_mul_5_p <= Pix_144;
    10'd5:  neuron_1_mul_5_p <= Pix_145;
    10'd6:  neuron_1_mul_5_p <= Pix_146;
    10'd7:  neuron_1_mul_5_p <= Pix_147;
    10'd8:  neuron_1_mul_5_p <= Pix_148;
    10'd9:  neuron_1_mul_5_p <= Pix_149;
    10'd10:  neuron_1_mul_5_p <= Pix_150;
    10'd11:  neuron_1_mul_5_p <= Pix_151;
    10'd12:  neuron_1_mul_5_p <= Pix_152;
    10'd13:  neuron_1_mul_5_p <= Pix_153;
    10'd14:  neuron_1_mul_5_p <= Pix_154;
    10'd15:  neuron_1_mul_5_p <= Pix_155;
    10'd16:  neuron_1_mul_5_p <= Pix_156;
    10'd17:  neuron_1_mul_5_p <= Pix_157;
    10'd18:  neuron_1_mul_5_p <= Pix_158;
    10'd19:  neuron_1_mul_5_p <= Pix_159;
    10'd20:  neuron_1_mul_5_p <= Pix_160;
    10'd21:  neuron_1_mul_5_p <= Pix_161;
    10'd22:  neuron_1_mul_5_p <= Pix_162;
    10'd23:  neuron_1_mul_5_p <= Pix_163;
    10'd24:  neuron_1_mul_5_p <= Pix_164;
    10'd25:  neuron_1_mul_5_p <= Pix_165;
    10'd26:  neuron_1_mul_5_p <= Pix_166;
    10'd27:  neuron_1_mul_5_p <= Pix_167;
    default: neuron_1_mul_5_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_6_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_6_p <= Pix_168;
    10'd1:  neuron_1_mul_6_p <= Pix_169;
    10'd2:  neuron_1_mul_6_p <= Pix_170;
    10'd3:  neuron_1_mul_6_p <= Pix_171;
    10'd4:  neuron_1_mul_6_p <= Pix_172;
    10'd5:  neuron_1_mul_6_p <= Pix_173;
    10'd6:  neuron_1_mul_6_p <= Pix_174;
    10'd7:  neuron_1_mul_6_p <= Pix_175;
    10'd8:  neuron_1_mul_6_p <= Pix_176;
    10'd9:  neuron_1_mul_6_p <= Pix_177;
    10'd10:  neuron_1_mul_6_p <= Pix_178;
    10'd11:  neuron_1_mul_6_p <= Pix_179;
    10'd12:  neuron_1_mul_6_p <= Pix_180;
    10'd13:  neuron_1_mul_6_p <= Pix_181;
    10'd14:  neuron_1_mul_6_p <= Pix_182;
    10'd15:  neuron_1_mul_6_p <= Pix_183;
    10'd16:  neuron_1_mul_6_p <= Pix_184;
    10'd17:  neuron_1_mul_6_p <= Pix_185;
    10'd18:  neuron_1_mul_6_p <= Pix_186;
    10'd19:  neuron_1_mul_6_p <= Pix_187;
    10'd20:  neuron_1_mul_6_p <= Pix_188;
    10'd21:  neuron_1_mul_6_p <= Pix_189;
    10'd22:  neuron_1_mul_6_p <= Pix_190;
    10'd23:  neuron_1_mul_6_p <= Pix_191;
    10'd24:  neuron_1_mul_6_p <= Pix_192;
    10'd25:  neuron_1_mul_6_p <= Pix_193;
    10'd26:  neuron_1_mul_6_p <= Pix_194;
    10'd27:  neuron_1_mul_6_p <= Pix_195;
    default: neuron_1_mul_6_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_7_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_7_p <= Pix_196;
    10'd1:  neuron_1_mul_7_p <= Pix_197;
    10'd2:  neuron_1_mul_7_p <= Pix_198;
    10'd3:  neuron_1_mul_7_p <= Pix_199;
    10'd4:  neuron_1_mul_7_p <= Pix_200;
    10'd5:  neuron_1_mul_7_p <= Pix_201;
    10'd6:  neuron_1_mul_7_p <= Pix_202;
    10'd7:  neuron_1_mul_7_p <= Pix_203;
    10'd8:  neuron_1_mul_7_p <= Pix_204;
    10'd9:  neuron_1_mul_7_p <= Pix_205;
    10'd10:  neuron_1_mul_7_p <= Pix_206;
    10'd11:  neuron_1_mul_7_p <= Pix_207;
    10'd12:  neuron_1_mul_7_p <= Pix_208;
    10'd13:  neuron_1_mul_7_p <= Pix_209;
    10'd14:  neuron_1_mul_7_p <= Pix_210;
    10'd15:  neuron_1_mul_7_p <= Pix_211;
    10'd16:  neuron_1_mul_7_p <= Pix_212;
    10'd17:  neuron_1_mul_7_p <= Pix_213;
    10'd18:  neuron_1_mul_7_p <= Pix_214;
    10'd19:  neuron_1_mul_7_p <= Pix_215;
    10'd20:  neuron_1_mul_7_p <= Pix_216;
    10'd21:  neuron_1_mul_7_p <= Pix_217;
    10'd22:  neuron_1_mul_7_p <= Pix_218;
    10'd23:  neuron_1_mul_7_p <= Pix_219;
    10'd24:  neuron_1_mul_7_p <= Pix_220;
    10'd25:  neuron_1_mul_7_p <= Pix_221;
    10'd26:  neuron_1_mul_7_p <= Pix_222;
    10'd27:  neuron_1_mul_7_p <= Pix_223;
    default: neuron_1_mul_7_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_8_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_8_p <= Pix_224;
    10'd1:  neuron_1_mul_8_p <= Pix_225;
    10'd2:  neuron_1_mul_8_p <= Pix_226;
    10'd3:  neuron_1_mul_8_p <= Pix_227;
    10'd4:  neuron_1_mul_8_p <= Pix_228;
    10'd5:  neuron_1_mul_8_p <= Pix_229;
    10'd6:  neuron_1_mul_8_p <= Pix_230;
    10'd7:  neuron_1_mul_8_p <= Pix_231;
    10'd8:  neuron_1_mul_8_p <= Pix_232;
    10'd9:  neuron_1_mul_8_p <= Pix_233;
    10'd10:  neuron_1_mul_8_p <= Pix_234;
    10'd11:  neuron_1_mul_8_p <= Pix_235;
    10'd12:  neuron_1_mul_8_p <= Pix_236;
    10'd13:  neuron_1_mul_8_p <= Pix_237;
    10'd14:  neuron_1_mul_8_p <= Pix_238;
    10'd15:  neuron_1_mul_8_p <= Pix_239;
    10'd16:  neuron_1_mul_8_p <= Pix_240;
    10'd17:  neuron_1_mul_8_p <= Pix_241;
    10'd18:  neuron_1_mul_8_p <= Pix_242;
    10'd19:  neuron_1_mul_8_p <= Pix_243;
    10'd20:  neuron_1_mul_8_p <= Pix_244;
    10'd21:  neuron_1_mul_8_p <= Pix_245;
    10'd22:  neuron_1_mul_8_p <= Pix_246;
    10'd23:  neuron_1_mul_8_p <= Pix_247;
    10'd24:  neuron_1_mul_8_p <= Pix_248;
    10'd25:  neuron_1_mul_8_p <= Pix_249;
    10'd26:  neuron_1_mul_8_p <= Pix_250;
    10'd27:  neuron_1_mul_8_p <= Pix_251;
    default: neuron_1_mul_8_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_9_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_9_p <= Pix_252;
    10'd1:  neuron_1_mul_9_p <= Pix_253;
    10'd2:  neuron_1_mul_9_p <= Pix_254;
    10'd3:  neuron_1_mul_9_p <= Pix_255;
    10'd4:  neuron_1_mul_9_p <= Pix_256;
    10'd5:  neuron_1_mul_9_p <= Pix_257;
    10'd6:  neuron_1_mul_9_p <= Pix_258;
    10'd7:  neuron_1_mul_9_p <= Pix_259;
    10'd8:  neuron_1_mul_9_p <= Pix_260;
    10'd9:  neuron_1_mul_9_p <= Pix_261;
    10'd10:  neuron_1_mul_9_p <= Pix_262;
    10'd11:  neuron_1_mul_9_p <= Pix_263;
    10'd12:  neuron_1_mul_9_p <= Pix_264;
    10'd13:  neuron_1_mul_9_p <= Pix_265;
    10'd14:  neuron_1_mul_9_p <= Pix_266;
    10'd15:  neuron_1_mul_9_p <= Pix_267;
    10'd16:  neuron_1_mul_9_p <= Pix_268;
    10'd17:  neuron_1_mul_9_p <= Pix_269;
    10'd18:  neuron_1_mul_9_p <= Pix_270;
    10'd19:  neuron_1_mul_9_p <= Pix_271;
    10'd20:  neuron_1_mul_9_p <= Pix_272;
    10'd21:  neuron_1_mul_9_p <= Pix_273;
    10'd22:  neuron_1_mul_9_p <= Pix_274;
    10'd23:  neuron_1_mul_9_p <= Pix_275;
    10'd24:  neuron_1_mul_9_p <= Pix_276;
    10'd25:  neuron_1_mul_9_p <= Pix_277;
    10'd26:  neuron_1_mul_9_p <= Pix_278;
    10'd27:  neuron_1_mul_9_p <= Pix_279;
    default: neuron_1_mul_9_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_10_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_10_p <= Pix_280;
    10'd1:  neuron_1_mul_10_p <= Pix_281;
    10'd2:  neuron_1_mul_10_p <= Pix_282;
    10'd3:  neuron_1_mul_10_p <= Pix_283;
    10'd4:  neuron_1_mul_10_p <= Pix_284;
    10'd5:  neuron_1_mul_10_p <= Pix_285;
    10'd6:  neuron_1_mul_10_p <= Pix_286;
    10'd7:  neuron_1_mul_10_p <= Pix_287;
    10'd8:  neuron_1_mul_10_p <= Pix_288;
    10'd9:  neuron_1_mul_10_p <= Pix_289;
    10'd10:  neuron_1_mul_10_p <= Pix_290;
    10'd11:  neuron_1_mul_10_p <= Pix_291;
    10'd12:  neuron_1_mul_10_p <= Pix_292;
    10'd13:  neuron_1_mul_10_p <= Pix_293;
    10'd14:  neuron_1_mul_10_p <= Pix_294;
    10'd15:  neuron_1_mul_10_p <= Pix_295;
    10'd16:  neuron_1_mul_10_p <= Pix_296;
    10'd17:  neuron_1_mul_10_p <= Pix_297;
    10'd18:  neuron_1_mul_10_p <= Pix_298;
    10'd19:  neuron_1_mul_10_p <= Pix_299;
    10'd20:  neuron_1_mul_10_p <= Pix_300;
    10'd21:  neuron_1_mul_10_p <= Pix_301;
    10'd22:  neuron_1_mul_10_p <= Pix_302;
    10'd23:  neuron_1_mul_10_p <= Pix_303;
    10'd24:  neuron_1_mul_10_p <= Pix_304;
    10'd25:  neuron_1_mul_10_p <= Pix_305;
    10'd26:  neuron_1_mul_10_p <= Pix_306;
    10'd27:  neuron_1_mul_10_p <= Pix_307;
    default: neuron_1_mul_10_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_11_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_11_p <= Pix_308;
    10'd1:  neuron_1_mul_11_p <= Pix_309;
    10'd2:  neuron_1_mul_11_p <= Pix_310;
    10'd3:  neuron_1_mul_11_p <= Pix_311;
    10'd4:  neuron_1_mul_11_p <= Pix_312;
    10'd5:  neuron_1_mul_11_p <= Pix_313;
    10'd6:  neuron_1_mul_11_p <= Pix_314;
    10'd7:  neuron_1_mul_11_p <= Pix_315;
    10'd8:  neuron_1_mul_11_p <= Pix_316;
    10'd9:  neuron_1_mul_11_p <= Pix_317;
    10'd10:  neuron_1_mul_11_p <= Pix_318;
    10'd11:  neuron_1_mul_11_p <= Pix_319;
    10'd12:  neuron_1_mul_11_p <= Pix_320;
    10'd13:  neuron_1_mul_11_p <= Pix_321;
    10'd14:  neuron_1_mul_11_p <= Pix_322;
    10'd15:  neuron_1_mul_11_p <= Pix_323;
    10'd16:  neuron_1_mul_11_p <= Pix_324;
    10'd17:  neuron_1_mul_11_p <= Pix_325;
    10'd18:  neuron_1_mul_11_p <= Pix_326;
    10'd19:  neuron_1_mul_11_p <= Pix_327;
    10'd20:  neuron_1_mul_11_p <= Pix_328;
    10'd21:  neuron_1_mul_11_p <= Pix_329;
    10'd22:  neuron_1_mul_11_p <= Pix_330;
    10'd23:  neuron_1_mul_11_p <= Pix_331;
    10'd24:  neuron_1_mul_11_p <= Pix_332;
    10'd25:  neuron_1_mul_11_p <= Pix_333;
    10'd26:  neuron_1_mul_11_p <= Pix_334;
    10'd27:  neuron_1_mul_11_p <= Pix_335;
    default: neuron_1_mul_11_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_12_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_12_p <= Pix_336;
    10'd1:  neuron_1_mul_12_p <= Pix_337;
    10'd2:  neuron_1_mul_12_p <= Pix_338;
    10'd3:  neuron_1_mul_12_p <= Pix_339;
    10'd4:  neuron_1_mul_12_p <= Pix_340;
    10'd5:  neuron_1_mul_12_p <= Pix_341;
    10'd6:  neuron_1_mul_12_p <= Pix_342;
    10'd7:  neuron_1_mul_12_p <= Pix_343;
    10'd8:  neuron_1_mul_12_p <= Pix_344;
    10'd9:  neuron_1_mul_12_p <= Pix_345;
    10'd10:  neuron_1_mul_12_p <= Pix_346;
    10'd11:  neuron_1_mul_12_p <= Pix_347;
    10'd12:  neuron_1_mul_12_p <= Pix_348;
    10'd13:  neuron_1_mul_12_p <= Pix_349;
    10'd14:  neuron_1_mul_12_p <= Pix_350;
    10'd15:  neuron_1_mul_12_p <= Pix_351;
    10'd16:  neuron_1_mul_12_p <= Pix_352;
    10'd17:  neuron_1_mul_12_p <= Pix_353;
    10'd18:  neuron_1_mul_12_p <= Pix_354;
    10'd19:  neuron_1_mul_12_p <= Pix_355;
    10'd20:  neuron_1_mul_12_p <= Pix_356;
    10'd21:  neuron_1_mul_12_p <= Pix_357;
    10'd22:  neuron_1_mul_12_p <= Pix_358;
    10'd23:  neuron_1_mul_12_p <= Pix_359;
    10'd24:  neuron_1_mul_12_p <= Pix_360;
    10'd25:  neuron_1_mul_12_p <= Pix_361;
    10'd26:  neuron_1_mul_12_p <= Pix_362;
    10'd27:  neuron_1_mul_12_p <= Pix_363;
    default: neuron_1_mul_12_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_13_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_13_p <= Pix_364;
    10'd1:  neuron_1_mul_13_p <= Pix_365;
    10'd2:  neuron_1_mul_13_p <= Pix_366;
    10'd3:  neuron_1_mul_13_p <= Pix_367;
    10'd4:  neuron_1_mul_13_p <= Pix_368;
    10'd5:  neuron_1_mul_13_p <= Pix_369;
    10'd6:  neuron_1_mul_13_p <= Pix_370;
    10'd7:  neuron_1_mul_13_p <= Pix_371;
    10'd8:  neuron_1_mul_13_p <= Pix_372;
    10'd9:  neuron_1_mul_13_p <= Pix_373;
    10'd10:  neuron_1_mul_13_p <= Pix_374;
    10'd11:  neuron_1_mul_13_p <= Pix_375;
    10'd12:  neuron_1_mul_13_p <= Pix_376;
    10'd13:  neuron_1_mul_13_p <= Pix_377;
    10'd14:  neuron_1_mul_13_p <= Pix_378;
    10'd15:  neuron_1_mul_13_p <= Pix_379;
    10'd16:  neuron_1_mul_13_p <= Pix_380;
    10'd17:  neuron_1_mul_13_p <= Pix_381;
    10'd18:  neuron_1_mul_13_p <= Pix_382;
    10'd19:  neuron_1_mul_13_p <= Pix_383;
    10'd20:  neuron_1_mul_13_p <= Pix_384;
    10'd21:  neuron_1_mul_13_p <= Pix_385;
    10'd22:  neuron_1_mul_13_p <= Pix_386;
    10'd23:  neuron_1_mul_13_p <= Pix_387;
    10'd24:  neuron_1_mul_13_p <= Pix_388;
    10'd25:  neuron_1_mul_13_p <= Pix_389;
    10'd26:  neuron_1_mul_13_p <= Pix_390;
    10'd27:  neuron_1_mul_13_p <= Pix_391;
    default: neuron_1_mul_13_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_14_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_14_p <= Pix_392;
    10'd1:  neuron_1_mul_14_p <= Pix_393;
    10'd2:  neuron_1_mul_14_p <= Pix_394;
    10'd3:  neuron_1_mul_14_p <= Pix_395;
    10'd4:  neuron_1_mul_14_p <= Pix_396;
    10'd5:  neuron_1_mul_14_p <= Pix_397;
    10'd6:  neuron_1_mul_14_p <= Pix_398;
    10'd7:  neuron_1_mul_14_p <= Pix_399;
    10'd8:  neuron_1_mul_14_p <= Pix_400;
    10'd9:  neuron_1_mul_14_p <= Pix_401;
    10'd10:  neuron_1_mul_14_p <= Pix_402;
    10'd11:  neuron_1_mul_14_p <= Pix_403;
    10'd12:  neuron_1_mul_14_p <= Pix_404;
    10'd13:  neuron_1_mul_14_p <= Pix_405;
    10'd14:  neuron_1_mul_14_p <= Pix_406;
    10'd15:  neuron_1_mul_14_p <= Pix_407;
    10'd16:  neuron_1_mul_14_p <= Pix_408;
    10'd17:  neuron_1_mul_14_p <= Pix_409;
    10'd18:  neuron_1_mul_14_p <= Pix_410;
    10'd19:  neuron_1_mul_14_p <= Pix_411;
    10'd20:  neuron_1_mul_14_p <= Pix_412;
    10'd21:  neuron_1_mul_14_p <= Pix_413;
    10'd22:  neuron_1_mul_14_p <= Pix_414;
    10'd23:  neuron_1_mul_14_p <= Pix_415;
    10'd24:  neuron_1_mul_14_p <= Pix_416;
    10'd25:  neuron_1_mul_14_p <= Pix_417;
    10'd26:  neuron_1_mul_14_p <= Pix_418;
    10'd27:  neuron_1_mul_14_p <= Pix_419;
    default: neuron_1_mul_14_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_15_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_15_p <= Pix_420;
    10'd1:  neuron_1_mul_15_p <= Pix_421;
    10'd2:  neuron_1_mul_15_p <= Pix_422;
    10'd3:  neuron_1_mul_15_p <= Pix_423;
    10'd4:  neuron_1_mul_15_p <= Pix_424;
    10'd5:  neuron_1_mul_15_p <= Pix_425;
    10'd6:  neuron_1_mul_15_p <= Pix_426;
    10'd7:  neuron_1_mul_15_p <= Pix_427;
    10'd8:  neuron_1_mul_15_p <= Pix_428;
    10'd9:  neuron_1_mul_15_p <= Pix_429;
    10'd10:  neuron_1_mul_15_p <= Pix_430;
    10'd11:  neuron_1_mul_15_p <= Pix_431;
    10'd12:  neuron_1_mul_15_p <= Pix_432;
    10'd13:  neuron_1_mul_15_p <= Pix_433;
    10'd14:  neuron_1_mul_15_p <= Pix_434;
    10'd15:  neuron_1_mul_15_p <= Pix_435;
    10'd16:  neuron_1_mul_15_p <= Pix_436;
    10'd17:  neuron_1_mul_15_p <= Pix_437;
    10'd18:  neuron_1_mul_15_p <= Pix_438;
    10'd19:  neuron_1_mul_15_p <= Pix_439;
    10'd20:  neuron_1_mul_15_p <= Pix_440;
    10'd21:  neuron_1_mul_15_p <= Pix_441;
    10'd22:  neuron_1_mul_15_p <= Pix_442;
    10'd23:  neuron_1_mul_15_p <= Pix_443;
    10'd24:  neuron_1_mul_15_p <= Pix_444;
    10'd25:  neuron_1_mul_15_p <= Pix_445;
    10'd26:  neuron_1_mul_15_p <= Pix_446;
    10'd27:  neuron_1_mul_15_p <= Pix_447;
    default: neuron_1_mul_15_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_16_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_16_p <= Pix_448;
    10'd1:  neuron_1_mul_16_p <= Pix_449;
    10'd2:  neuron_1_mul_16_p <= Pix_450;
    10'd3:  neuron_1_mul_16_p <= Pix_451;
    10'd4:  neuron_1_mul_16_p <= Pix_452;
    10'd5:  neuron_1_mul_16_p <= Pix_453;
    10'd6:  neuron_1_mul_16_p <= Pix_454;
    10'd7:  neuron_1_mul_16_p <= Pix_455;
    10'd8:  neuron_1_mul_16_p <= Pix_456;
    10'd9:  neuron_1_mul_16_p <= Pix_457;
    10'd10:  neuron_1_mul_16_p <= Pix_458;
    10'd11:  neuron_1_mul_16_p <= Pix_459;
    10'd12:  neuron_1_mul_16_p <= Pix_460;
    10'd13:  neuron_1_mul_16_p <= Pix_461;
    10'd14:  neuron_1_mul_16_p <= Pix_462;
    10'd15:  neuron_1_mul_16_p <= Pix_463;
    10'd16:  neuron_1_mul_16_p <= Pix_464;
    10'd17:  neuron_1_mul_16_p <= Pix_465;
    10'd18:  neuron_1_mul_16_p <= Pix_466;
    10'd19:  neuron_1_mul_16_p <= Pix_467;
    10'd20:  neuron_1_mul_16_p <= Pix_468;
    10'd21:  neuron_1_mul_16_p <= Pix_469;
    10'd22:  neuron_1_mul_16_p <= Pix_470;
    10'd23:  neuron_1_mul_16_p <= Pix_471;
    10'd24:  neuron_1_mul_16_p <= Pix_472;
    10'd25:  neuron_1_mul_16_p <= Pix_473;
    10'd26:  neuron_1_mul_16_p <= Pix_474;
    10'd27:  neuron_1_mul_16_p <= Pix_475;
    default: neuron_1_mul_16_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_17_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_17_p <= Pix_476;
    10'd1:  neuron_1_mul_17_p <= Pix_477;
    10'd2:  neuron_1_mul_17_p <= Pix_478;
    10'd3:  neuron_1_mul_17_p <= Pix_479;
    10'd4:  neuron_1_mul_17_p <= Pix_480;
    10'd5:  neuron_1_mul_17_p <= Pix_481;
    10'd6:  neuron_1_mul_17_p <= Pix_482;
    10'd7:  neuron_1_mul_17_p <= Pix_483;
    10'd8:  neuron_1_mul_17_p <= Pix_484;
    10'd9:  neuron_1_mul_17_p <= Pix_485;
    10'd10:  neuron_1_mul_17_p <= Pix_486;
    10'd11:  neuron_1_mul_17_p <= Pix_487;
    10'd12:  neuron_1_mul_17_p <= Pix_488;
    10'd13:  neuron_1_mul_17_p <= Pix_489;
    10'd14:  neuron_1_mul_17_p <= Pix_490;
    10'd15:  neuron_1_mul_17_p <= Pix_491;
    10'd16:  neuron_1_mul_17_p <= Pix_492;
    10'd17:  neuron_1_mul_17_p <= Pix_493;
    10'd18:  neuron_1_mul_17_p <= Pix_494;
    10'd19:  neuron_1_mul_17_p <= Pix_495;
    10'd20:  neuron_1_mul_17_p <= Pix_496;
    10'd21:  neuron_1_mul_17_p <= Pix_497;
    10'd22:  neuron_1_mul_17_p <= Pix_498;
    10'd23:  neuron_1_mul_17_p <= Pix_499;
    10'd24:  neuron_1_mul_17_p <= Pix_500;
    10'd25:  neuron_1_mul_17_p <= Pix_501;
    10'd26:  neuron_1_mul_17_p <= Pix_502;
    10'd27:  neuron_1_mul_17_p <= Pix_503;
    default: neuron_1_mul_17_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_18_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_18_p <= Pix_504;
    10'd1:  neuron_1_mul_18_p <= Pix_505;
    10'd2:  neuron_1_mul_18_p <= Pix_506;
    10'd3:  neuron_1_mul_18_p <= Pix_507;
    10'd4:  neuron_1_mul_18_p <= Pix_508;
    10'd5:  neuron_1_mul_18_p <= Pix_509;
    10'd6:  neuron_1_mul_18_p <= Pix_510;
    10'd7:  neuron_1_mul_18_p <= Pix_511;
    10'd8:  neuron_1_mul_18_p <= Pix_512;
    10'd9:  neuron_1_mul_18_p <= Pix_513;
    10'd10:  neuron_1_mul_18_p <= Pix_514;
    10'd11:  neuron_1_mul_18_p <= Pix_515;
    10'd12:  neuron_1_mul_18_p <= Pix_516;
    10'd13:  neuron_1_mul_18_p <= Pix_517;
    10'd14:  neuron_1_mul_18_p <= Pix_518;
    10'd15:  neuron_1_mul_18_p <= Pix_519;
    10'd16:  neuron_1_mul_18_p <= Pix_520;
    10'd17:  neuron_1_mul_18_p <= Pix_521;
    10'd18:  neuron_1_mul_18_p <= Pix_522;
    10'd19:  neuron_1_mul_18_p <= Pix_523;
    10'd20:  neuron_1_mul_18_p <= Pix_524;
    10'd21:  neuron_1_mul_18_p <= Pix_525;
    10'd22:  neuron_1_mul_18_p <= Pix_526;
    10'd23:  neuron_1_mul_18_p <= Pix_527;
    10'd24:  neuron_1_mul_18_p <= Pix_528;
    10'd25:  neuron_1_mul_18_p <= Pix_529;
    10'd26:  neuron_1_mul_18_p <= Pix_530;
    10'd27:  neuron_1_mul_18_p <= Pix_531;
    default: neuron_1_mul_18_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_19_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_19_p <= Pix_532;
    10'd1:  neuron_1_mul_19_p <= Pix_533;
    10'd2:  neuron_1_mul_19_p <= Pix_534;
    10'd3:  neuron_1_mul_19_p <= Pix_535;
    10'd4:  neuron_1_mul_19_p <= Pix_536;
    10'd5:  neuron_1_mul_19_p <= Pix_537;
    10'd6:  neuron_1_mul_19_p <= Pix_538;
    10'd7:  neuron_1_mul_19_p <= Pix_539;
    10'd8:  neuron_1_mul_19_p <= Pix_540;
    10'd9:  neuron_1_mul_19_p <= Pix_541;
    10'd10:  neuron_1_mul_19_p <= Pix_542;
    10'd11:  neuron_1_mul_19_p <= Pix_543;
    10'd12:  neuron_1_mul_19_p <= Pix_544;
    10'd13:  neuron_1_mul_19_p <= Pix_545;
    10'd14:  neuron_1_mul_19_p <= Pix_546;
    10'd15:  neuron_1_mul_19_p <= Pix_547;
    10'd16:  neuron_1_mul_19_p <= Pix_548;
    10'd17:  neuron_1_mul_19_p <= Pix_549;
    10'd18:  neuron_1_mul_19_p <= Pix_550;
    10'd19:  neuron_1_mul_19_p <= Pix_551;
    10'd20:  neuron_1_mul_19_p <= Pix_552;
    10'd21:  neuron_1_mul_19_p <= Pix_553;
    10'd22:  neuron_1_mul_19_p <= Pix_554;
    10'd23:  neuron_1_mul_19_p <= Pix_555;
    10'd24:  neuron_1_mul_19_p <= Pix_556;
    10'd25:  neuron_1_mul_19_p <= Pix_557;
    10'd26:  neuron_1_mul_19_p <= Pix_558;
    10'd27:  neuron_1_mul_19_p <= Pix_559;
    default: neuron_1_mul_19_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_20_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_20_p <= Pix_560;
    10'd1:  neuron_1_mul_20_p <= Pix_561;
    10'd2:  neuron_1_mul_20_p <= Pix_562;
    10'd3:  neuron_1_mul_20_p <= Pix_563;
    10'd4:  neuron_1_mul_20_p <= Pix_564;
    10'd5:  neuron_1_mul_20_p <= Pix_565;
    10'd6:  neuron_1_mul_20_p <= Pix_566;
    10'd7:  neuron_1_mul_20_p <= Pix_567;
    10'd8:  neuron_1_mul_20_p <= Pix_568;
    10'd9:  neuron_1_mul_20_p <= Pix_569;
    10'd10:  neuron_1_mul_20_p <= Pix_570;
    10'd11:  neuron_1_mul_20_p <= Pix_571;
    10'd12:  neuron_1_mul_20_p <= Pix_572;
    10'd13:  neuron_1_mul_20_p <= Pix_573;
    10'd14:  neuron_1_mul_20_p <= Pix_574;
    10'd15:  neuron_1_mul_20_p <= Pix_575;
    10'd16:  neuron_1_mul_20_p <= Pix_576;
    10'd17:  neuron_1_mul_20_p <= Pix_577;
    10'd18:  neuron_1_mul_20_p <= Pix_578;
    10'd19:  neuron_1_mul_20_p <= Pix_579;
    10'd20:  neuron_1_mul_20_p <= Pix_580;
    10'd21:  neuron_1_mul_20_p <= Pix_581;
    10'd22:  neuron_1_mul_20_p <= Pix_582;
    10'd23:  neuron_1_mul_20_p <= Pix_583;
    10'd24:  neuron_1_mul_20_p <= Pix_584;
    10'd25:  neuron_1_mul_20_p <= Pix_585;
    10'd26:  neuron_1_mul_20_p <= Pix_586;
    10'd27:  neuron_1_mul_20_p <= Pix_587;
    default: neuron_1_mul_20_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_21_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_21_p <= Pix_588;
    10'd1:  neuron_1_mul_21_p <= Pix_589;
    10'd2:  neuron_1_mul_21_p <= Pix_590;
    10'd3:  neuron_1_mul_21_p <= Pix_591;
    10'd4:  neuron_1_mul_21_p <= Pix_592;
    10'd5:  neuron_1_mul_21_p <= Pix_593;
    10'd6:  neuron_1_mul_21_p <= Pix_594;
    10'd7:  neuron_1_mul_21_p <= Pix_595;
    10'd8:  neuron_1_mul_21_p <= Pix_596;
    10'd9:  neuron_1_mul_21_p <= Pix_597;
    10'd10:  neuron_1_mul_21_p <= Pix_598;
    10'd11:  neuron_1_mul_21_p <= Pix_599;
    10'd12:  neuron_1_mul_21_p <= Pix_600;
    10'd13:  neuron_1_mul_21_p <= Pix_601;
    10'd14:  neuron_1_mul_21_p <= Pix_602;
    10'd15:  neuron_1_mul_21_p <= Pix_603;
    10'd16:  neuron_1_mul_21_p <= Pix_604;
    10'd17:  neuron_1_mul_21_p <= Pix_605;
    10'd18:  neuron_1_mul_21_p <= Pix_606;
    10'd19:  neuron_1_mul_21_p <= Pix_607;
    10'd20:  neuron_1_mul_21_p <= Pix_608;
    10'd21:  neuron_1_mul_21_p <= Pix_609;
    10'd22:  neuron_1_mul_21_p <= Pix_610;
    10'd23:  neuron_1_mul_21_p <= Pix_611;
    10'd24:  neuron_1_mul_21_p <= Pix_612;
    10'd25:  neuron_1_mul_21_p <= Pix_613;
    10'd26:  neuron_1_mul_21_p <= Pix_614;
    10'd27:  neuron_1_mul_21_p <= Pix_615;
    default: neuron_1_mul_21_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_22_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_22_p <= Pix_616;
    10'd1:  neuron_1_mul_22_p <= Pix_617;
    10'd2:  neuron_1_mul_22_p <= Pix_618;
    10'd3:  neuron_1_mul_22_p <= Pix_619;
    10'd4:  neuron_1_mul_22_p <= Pix_620;
    10'd5:  neuron_1_mul_22_p <= Pix_621;
    10'd6:  neuron_1_mul_22_p <= Pix_622;
    10'd7:  neuron_1_mul_22_p <= Pix_623;
    10'd8:  neuron_1_mul_22_p <= Pix_624;
    10'd9:  neuron_1_mul_22_p <= Pix_625;
    10'd10:  neuron_1_mul_22_p <= Pix_626;
    10'd11:  neuron_1_mul_22_p <= Pix_627;
    10'd12:  neuron_1_mul_22_p <= Pix_628;
    10'd13:  neuron_1_mul_22_p <= Pix_629;
    10'd14:  neuron_1_mul_22_p <= Pix_630;
    10'd15:  neuron_1_mul_22_p <= Pix_631;
    10'd16:  neuron_1_mul_22_p <= Pix_632;
    10'd17:  neuron_1_mul_22_p <= Pix_633;
    10'd18:  neuron_1_mul_22_p <= Pix_634;
    10'd19:  neuron_1_mul_22_p <= Pix_635;
    10'd20:  neuron_1_mul_22_p <= Pix_636;
    10'd21:  neuron_1_mul_22_p <= Pix_637;
    10'd22:  neuron_1_mul_22_p <= Pix_638;
    10'd23:  neuron_1_mul_22_p <= Pix_639;
    10'd24:  neuron_1_mul_22_p <= Pix_640;
    10'd25:  neuron_1_mul_22_p <= Pix_641;
    10'd26:  neuron_1_mul_22_p <= Pix_642;
    10'd27:  neuron_1_mul_22_p <= Pix_643;
    default: neuron_1_mul_22_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_23_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_23_p <= Pix_644;
    10'd1:  neuron_1_mul_23_p <= Pix_645;
    10'd2:  neuron_1_mul_23_p <= Pix_646;
    10'd3:  neuron_1_mul_23_p <= Pix_647;
    10'd4:  neuron_1_mul_23_p <= Pix_648;
    10'd5:  neuron_1_mul_23_p <= Pix_649;
    10'd6:  neuron_1_mul_23_p <= Pix_650;
    10'd7:  neuron_1_mul_23_p <= Pix_651;
    10'd8:  neuron_1_mul_23_p <= Pix_652;
    10'd9:  neuron_1_mul_23_p <= Pix_653;
    10'd10:  neuron_1_mul_23_p <= Pix_654;
    10'd11:  neuron_1_mul_23_p <= Pix_655;
    10'd12:  neuron_1_mul_23_p <= Pix_656;
    10'd13:  neuron_1_mul_23_p <= Pix_657;
    10'd14:  neuron_1_mul_23_p <= Pix_658;
    10'd15:  neuron_1_mul_23_p <= Pix_659;
    10'd16:  neuron_1_mul_23_p <= Pix_660;
    10'd17:  neuron_1_mul_23_p <= Pix_661;
    10'd18:  neuron_1_mul_23_p <= Pix_662;
    10'd19:  neuron_1_mul_23_p <= Pix_663;
    10'd20:  neuron_1_mul_23_p <= Pix_664;
    10'd21:  neuron_1_mul_23_p <= Pix_665;
    10'd22:  neuron_1_mul_23_p <= Pix_666;
    10'd23:  neuron_1_mul_23_p <= Pix_667;
    10'd24:  neuron_1_mul_23_p <= Pix_668;
    10'd25:  neuron_1_mul_23_p <= Pix_669;
    10'd26:  neuron_1_mul_23_p <= Pix_670;
    10'd27:  neuron_1_mul_23_p <= Pix_671;
    default: neuron_1_mul_23_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_24_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_24_p <= Pix_672;
    10'd1:  neuron_1_mul_24_p <= Pix_673;
    10'd2:  neuron_1_mul_24_p <= Pix_674;
    10'd3:  neuron_1_mul_24_p <= Pix_675;
    10'd4:  neuron_1_mul_24_p <= Pix_676;
    10'd5:  neuron_1_mul_24_p <= Pix_677;
    10'd6:  neuron_1_mul_24_p <= Pix_678;
    10'd7:  neuron_1_mul_24_p <= Pix_679;
    10'd8:  neuron_1_mul_24_p <= Pix_680;
    10'd9:  neuron_1_mul_24_p <= Pix_681;
    10'd10:  neuron_1_mul_24_p <= Pix_682;
    10'd11:  neuron_1_mul_24_p <= Pix_683;
    10'd12:  neuron_1_mul_24_p <= Pix_684;
    10'd13:  neuron_1_mul_24_p <= Pix_685;
    10'd14:  neuron_1_mul_24_p <= Pix_686;
    10'd15:  neuron_1_mul_24_p <= Pix_687;
    10'd16:  neuron_1_mul_24_p <= Pix_688;
    10'd17:  neuron_1_mul_24_p <= Pix_689;
    10'd18:  neuron_1_mul_24_p <= Pix_690;
    10'd19:  neuron_1_mul_24_p <= Pix_691;
    10'd20:  neuron_1_mul_24_p <= Pix_692;
    10'd21:  neuron_1_mul_24_p <= Pix_693;
    10'd22:  neuron_1_mul_24_p <= Pix_694;
    10'd23:  neuron_1_mul_24_p <= Pix_695;
    10'd24:  neuron_1_mul_24_p <= Pix_696;
    10'd25:  neuron_1_mul_24_p <= Pix_697;
    10'd26:  neuron_1_mul_24_p <= Pix_698;
    10'd27:  neuron_1_mul_24_p <= Pix_699;
    default: neuron_1_mul_24_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_25_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_25_p <= Pix_700;
    10'd1:  neuron_1_mul_25_p <= Pix_701;
    10'd2:  neuron_1_mul_25_p <= Pix_702;
    10'd3:  neuron_1_mul_25_p <= Pix_703;
    10'd4:  neuron_1_mul_25_p <= Pix_704;
    10'd5:  neuron_1_mul_25_p <= Pix_705;
    10'd6:  neuron_1_mul_25_p <= Pix_706;
    10'd7:  neuron_1_mul_25_p <= Pix_707;
    10'd8:  neuron_1_mul_25_p <= Pix_708;
    10'd9:  neuron_1_mul_25_p <= Pix_709;
    10'd10:  neuron_1_mul_25_p <= Pix_710;
    10'd11:  neuron_1_mul_25_p <= Pix_711;
    10'd12:  neuron_1_mul_25_p <= Pix_712;
    10'd13:  neuron_1_mul_25_p <= Pix_713;
    10'd14:  neuron_1_mul_25_p <= Pix_714;
    10'd15:  neuron_1_mul_25_p <= Pix_715;
    10'd16:  neuron_1_mul_25_p <= Pix_716;
    10'd17:  neuron_1_mul_25_p <= Pix_717;
    10'd18:  neuron_1_mul_25_p <= Pix_718;
    10'd19:  neuron_1_mul_25_p <= Pix_719;
    10'd20:  neuron_1_mul_25_p <= Pix_720;
    10'd21:  neuron_1_mul_25_p <= Pix_721;
    10'd22:  neuron_1_mul_25_p <= Pix_722;
    10'd23:  neuron_1_mul_25_p <= Pix_723;
    10'd24:  neuron_1_mul_25_p <= Pix_724;
    10'd25:  neuron_1_mul_25_p <= Pix_725;
    10'd26:  neuron_1_mul_25_p <= Pix_726;
    10'd27:  neuron_1_mul_25_p <= Pix_727;
    default: neuron_1_mul_25_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_26_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_26_p <= Pix_728;
    10'd1:  neuron_1_mul_26_p <= Pix_729;
    10'd2:  neuron_1_mul_26_p <= Pix_730;
    10'd3:  neuron_1_mul_26_p <= Pix_731;
    10'd4:  neuron_1_mul_26_p <= Pix_732;
    10'd5:  neuron_1_mul_26_p <= Pix_733;
    10'd6:  neuron_1_mul_26_p <= Pix_734;
    10'd7:  neuron_1_mul_26_p <= Pix_735;
    10'd8:  neuron_1_mul_26_p <= Pix_736;
    10'd9:  neuron_1_mul_26_p <= Pix_737;
    10'd10:  neuron_1_mul_26_p <= Pix_738;
    10'd11:  neuron_1_mul_26_p <= Pix_739;
    10'd12:  neuron_1_mul_26_p <= Pix_740;
    10'd13:  neuron_1_mul_26_p <= Pix_741;
    10'd14:  neuron_1_mul_26_p <= Pix_742;
    10'd15:  neuron_1_mul_26_p <= Pix_743;
    10'd16:  neuron_1_mul_26_p <= Pix_744;
    10'd17:  neuron_1_mul_26_p <= Pix_745;
    10'd18:  neuron_1_mul_26_p <= Pix_746;
    10'd19:  neuron_1_mul_26_p <= Pix_747;
    10'd20:  neuron_1_mul_26_p <= Pix_748;
    10'd21:  neuron_1_mul_26_p <= Pix_749;
    10'd22:  neuron_1_mul_26_p <= Pix_750;
    10'd23:  neuron_1_mul_26_p <= Pix_751;
    10'd24:  neuron_1_mul_26_p <= Pix_752;
    10'd25:  neuron_1_mul_26_p <= Pix_753;
    10'd26:  neuron_1_mul_26_p <= Pix_754;
    10'd27:  neuron_1_mul_26_p <= Pix_755;
    default: neuron_1_mul_26_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_1_mul_27_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_1_mul_27_p <= Pix_756;
    10'd1:  neuron_1_mul_27_p <= Pix_757;
    10'd2:  neuron_1_mul_27_p <= Pix_758;
    10'd3:  neuron_1_mul_27_p <= Pix_759;
    10'd4:  neuron_1_mul_27_p <= Pix_760;
    10'd5:  neuron_1_mul_27_p <= Pix_761;
    10'd6:  neuron_1_mul_27_p <= Pix_762;
    10'd7:  neuron_1_mul_27_p <= Pix_763;
    10'd8:  neuron_1_mul_27_p <= Pix_764;
    10'd9:  neuron_1_mul_27_p <= Pix_765;
    10'd10:  neuron_1_mul_27_p <= Pix_766;
    10'd11:  neuron_1_mul_27_p <= Pix_767;
    10'd12:  neuron_1_mul_27_p <= Pix_768;
    10'd13:  neuron_1_mul_27_p <= Pix_769;
    10'd14:  neuron_1_mul_27_p <= Pix_770;
    10'd15:  neuron_1_mul_27_p <= Pix_771;
    10'd16:  neuron_1_mul_27_p <= Pix_772;
    10'd17:  neuron_1_mul_27_p <= Pix_773;
    10'd18:  neuron_1_mul_27_p <= Pix_774;
    10'd19:  neuron_1_mul_27_p <= Pix_775;
    10'd20:  neuron_1_mul_27_p <= Pix_776;
    10'd21:  neuron_1_mul_27_p <= Pix_777;
    10'd22:  neuron_1_mul_27_p <= Pix_778;
    10'd23:  neuron_1_mul_27_p <= Pix_779;
    10'd24:  neuron_1_mul_27_p <= Pix_780;
    10'd25:  neuron_1_mul_27_p <= Pix_781;
    10'd26:  neuron_1_mul_27_p <= Pix_782;
    10'd27:  neuron_1_mul_27_p <= Pix_783;
    default: neuron_1_mul_27_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_0_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_0_p <= Pix_0;
    10'd1:  neuron_2_mul_0_p <= Pix_1;
    10'd2:  neuron_2_mul_0_p <= Pix_2;
    10'd3:  neuron_2_mul_0_p <= Pix_3;
    10'd4:  neuron_2_mul_0_p <= Pix_4;
    10'd5:  neuron_2_mul_0_p <= Pix_5;
    10'd6:  neuron_2_mul_0_p <= Pix_6;
    10'd7:  neuron_2_mul_0_p <= Pix_7;
    10'd8:  neuron_2_mul_0_p <= Pix_8;
    10'd9:  neuron_2_mul_0_p <= Pix_9;
    10'd10:  neuron_2_mul_0_p <= Pix_10;
    10'd11:  neuron_2_mul_0_p <= Pix_11;
    10'd12:  neuron_2_mul_0_p <= Pix_12;
    10'd13:  neuron_2_mul_0_p <= Pix_13;
    10'd14:  neuron_2_mul_0_p <= Pix_14;
    10'd15:  neuron_2_mul_0_p <= Pix_15;
    10'd16:  neuron_2_mul_0_p <= Pix_16;
    10'd17:  neuron_2_mul_0_p <= Pix_17;
    10'd18:  neuron_2_mul_0_p <= Pix_18;
    10'd19:  neuron_2_mul_0_p <= Pix_19;
    10'd20:  neuron_2_mul_0_p <= Pix_20;
    10'd21:  neuron_2_mul_0_p <= Pix_21;
    10'd22:  neuron_2_mul_0_p <= Pix_22;
    10'd23:  neuron_2_mul_0_p <= Pix_23;
    10'd24:  neuron_2_mul_0_p <= Pix_24;
    10'd25:  neuron_2_mul_0_p <= Pix_25;
    10'd26:  neuron_2_mul_0_p <= Pix_26;
    10'd27:  neuron_2_mul_0_p <= Pix_27;
    default: neuron_2_mul_0_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_1_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_1_p <= Pix_28;
    10'd1:  neuron_2_mul_1_p <= Pix_29;
    10'd2:  neuron_2_mul_1_p <= Pix_30;
    10'd3:  neuron_2_mul_1_p <= Pix_31;
    10'd4:  neuron_2_mul_1_p <= Pix_32;
    10'd5:  neuron_2_mul_1_p <= Pix_33;
    10'd6:  neuron_2_mul_1_p <= Pix_34;
    10'd7:  neuron_2_mul_1_p <= Pix_35;
    10'd8:  neuron_2_mul_1_p <= Pix_36;
    10'd9:  neuron_2_mul_1_p <= Pix_37;
    10'd10:  neuron_2_mul_1_p <= Pix_38;
    10'd11:  neuron_2_mul_1_p <= Pix_39;
    10'd12:  neuron_2_mul_1_p <= Pix_40;
    10'd13:  neuron_2_mul_1_p <= Pix_41;
    10'd14:  neuron_2_mul_1_p <= Pix_42;
    10'd15:  neuron_2_mul_1_p <= Pix_43;
    10'd16:  neuron_2_mul_1_p <= Pix_44;
    10'd17:  neuron_2_mul_1_p <= Pix_45;
    10'd18:  neuron_2_mul_1_p <= Pix_46;
    10'd19:  neuron_2_mul_1_p <= Pix_47;
    10'd20:  neuron_2_mul_1_p <= Pix_48;
    10'd21:  neuron_2_mul_1_p <= Pix_49;
    10'd22:  neuron_2_mul_1_p <= Pix_50;
    10'd23:  neuron_2_mul_1_p <= Pix_51;
    10'd24:  neuron_2_mul_1_p <= Pix_52;
    10'd25:  neuron_2_mul_1_p <= Pix_53;
    10'd26:  neuron_2_mul_1_p <= Pix_54;
    10'd27:  neuron_2_mul_1_p <= Pix_55;
    default: neuron_2_mul_1_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_2_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_2_p <= Pix_56;
    10'd1:  neuron_2_mul_2_p <= Pix_57;
    10'd2:  neuron_2_mul_2_p <= Pix_58;
    10'd3:  neuron_2_mul_2_p <= Pix_59;
    10'd4:  neuron_2_mul_2_p <= Pix_60;
    10'd5:  neuron_2_mul_2_p <= Pix_61;
    10'd6:  neuron_2_mul_2_p <= Pix_62;
    10'd7:  neuron_2_mul_2_p <= Pix_63;
    10'd8:  neuron_2_mul_2_p <= Pix_64;
    10'd9:  neuron_2_mul_2_p <= Pix_65;
    10'd10:  neuron_2_mul_2_p <= Pix_66;
    10'd11:  neuron_2_mul_2_p <= Pix_67;
    10'd12:  neuron_2_mul_2_p <= Pix_68;
    10'd13:  neuron_2_mul_2_p <= Pix_69;
    10'd14:  neuron_2_mul_2_p <= Pix_70;
    10'd15:  neuron_2_mul_2_p <= Pix_71;
    10'd16:  neuron_2_mul_2_p <= Pix_72;
    10'd17:  neuron_2_mul_2_p <= Pix_73;
    10'd18:  neuron_2_mul_2_p <= Pix_74;
    10'd19:  neuron_2_mul_2_p <= Pix_75;
    10'd20:  neuron_2_mul_2_p <= Pix_76;
    10'd21:  neuron_2_mul_2_p <= Pix_77;
    10'd22:  neuron_2_mul_2_p <= Pix_78;
    10'd23:  neuron_2_mul_2_p <= Pix_79;
    10'd24:  neuron_2_mul_2_p <= Pix_80;
    10'd25:  neuron_2_mul_2_p <= Pix_81;
    10'd26:  neuron_2_mul_2_p <= Pix_82;
    10'd27:  neuron_2_mul_2_p <= Pix_83;
    default: neuron_2_mul_2_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_3_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_3_p <= Pix_84;
    10'd1:  neuron_2_mul_3_p <= Pix_85;
    10'd2:  neuron_2_mul_3_p <= Pix_86;
    10'd3:  neuron_2_mul_3_p <= Pix_87;
    10'd4:  neuron_2_mul_3_p <= Pix_88;
    10'd5:  neuron_2_mul_3_p <= Pix_89;
    10'd6:  neuron_2_mul_3_p <= Pix_90;
    10'd7:  neuron_2_mul_3_p <= Pix_91;
    10'd8:  neuron_2_mul_3_p <= Pix_92;
    10'd9:  neuron_2_mul_3_p <= Pix_93;
    10'd10:  neuron_2_mul_3_p <= Pix_94;
    10'd11:  neuron_2_mul_3_p <= Pix_95;
    10'd12:  neuron_2_mul_3_p <= Pix_96;
    10'd13:  neuron_2_mul_3_p <= Pix_97;
    10'd14:  neuron_2_mul_3_p <= Pix_98;
    10'd15:  neuron_2_mul_3_p <= Pix_99;
    10'd16:  neuron_2_mul_3_p <= Pix_100;
    10'd17:  neuron_2_mul_3_p <= Pix_101;
    10'd18:  neuron_2_mul_3_p <= Pix_102;
    10'd19:  neuron_2_mul_3_p <= Pix_103;
    10'd20:  neuron_2_mul_3_p <= Pix_104;
    10'd21:  neuron_2_mul_3_p <= Pix_105;
    10'd22:  neuron_2_mul_3_p <= Pix_106;
    10'd23:  neuron_2_mul_3_p <= Pix_107;
    10'd24:  neuron_2_mul_3_p <= Pix_108;
    10'd25:  neuron_2_mul_3_p <= Pix_109;
    10'd26:  neuron_2_mul_3_p <= Pix_110;
    10'd27:  neuron_2_mul_3_p <= Pix_111;
    default: neuron_2_mul_3_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_4_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_4_p <= Pix_112;
    10'd1:  neuron_2_mul_4_p <= Pix_113;
    10'd2:  neuron_2_mul_4_p <= Pix_114;
    10'd3:  neuron_2_mul_4_p <= Pix_115;
    10'd4:  neuron_2_mul_4_p <= Pix_116;
    10'd5:  neuron_2_mul_4_p <= Pix_117;
    10'd6:  neuron_2_mul_4_p <= Pix_118;
    10'd7:  neuron_2_mul_4_p <= Pix_119;
    10'd8:  neuron_2_mul_4_p <= Pix_120;
    10'd9:  neuron_2_mul_4_p <= Pix_121;
    10'd10:  neuron_2_mul_4_p <= Pix_122;
    10'd11:  neuron_2_mul_4_p <= Pix_123;
    10'd12:  neuron_2_mul_4_p <= Pix_124;
    10'd13:  neuron_2_mul_4_p <= Pix_125;
    10'd14:  neuron_2_mul_4_p <= Pix_126;
    10'd15:  neuron_2_mul_4_p <= Pix_127;
    10'd16:  neuron_2_mul_4_p <= Pix_128;
    10'd17:  neuron_2_mul_4_p <= Pix_129;
    10'd18:  neuron_2_mul_4_p <= Pix_130;
    10'd19:  neuron_2_mul_4_p <= Pix_131;
    10'd20:  neuron_2_mul_4_p <= Pix_132;
    10'd21:  neuron_2_mul_4_p <= Pix_133;
    10'd22:  neuron_2_mul_4_p <= Pix_134;
    10'd23:  neuron_2_mul_4_p <= Pix_135;
    10'd24:  neuron_2_mul_4_p <= Pix_136;
    10'd25:  neuron_2_mul_4_p <= Pix_137;
    10'd26:  neuron_2_mul_4_p <= Pix_138;
    10'd27:  neuron_2_mul_4_p <= Pix_139;
    default: neuron_2_mul_4_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_5_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_5_p <= Pix_140;
    10'd1:  neuron_2_mul_5_p <= Pix_141;
    10'd2:  neuron_2_mul_5_p <= Pix_142;
    10'd3:  neuron_2_mul_5_p <= Pix_143;
    10'd4:  neuron_2_mul_5_p <= Pix_144;
    10'd5:  neuron_2_mul_5_p <= Pix_145;
    10'd6:  neuron_2_mul_5_p <= Pix_146;
    10'd7:  neuron_2_mul_5_p <= Pix_147;
    10'd8:  neuron_2_mul_5_p <= Pix_148;
    10'd9:  neuron_2_mul_5_p <= Pix_149;
    10'd10:  neuron_2_mul_5_p <= Pix_150;
    10'd11:  neuron_2_mul_5_p <= Pix_151;
    10'd12:  neuron_2_mul_5_p <= Pix_152;
    10'd13:  neuron_2_mul_5_p <= Pix_153;
    10'd14:  neuron_2_mul_5_p <= Pix_154;
    10'd15:  neuron_2_mul_5_p <= Pix_155;
    10'd16:  neuron_2_mul_5_p <= Pix_156;
    10'd17:  neuron_2_mul_5_p <= Pix_157;
    10'd18:  neuron_2_mul_5_p <= Pix_158;
    10'd19:  neuron_2_mul_5_p <= Pix_159;
    10'd20:  neuron_2_mul_5_p <= Pix_160;
    10'd21:  neuron_2_mul_5_p <= Pix_161;
    10'd22:  neuron_2_mul_5_p <= Pix_162;
    10'd23:  neuron_2_mul_5_p <= Pix_163;
    10'd24:  neuron_2_mul_5_p <= Pix_164;
    10'd25:  neuron_2_mul_5_p <= Pix_165;
    10'd26:  neuron_2_mul_5_p <= Pix_166;
    10'd27:  neuron_2_mul_5_p <= Pix_167;
    default: neuron_2_mul_5_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_6_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_6_p <= Pix_168;
    10'd1:  neuron_2_mul_6_p <= Pix_169;
    10'd2:  neuron_2_mul_6_p <= Pix_170;
    10'd3:  neuron_2_mul_6_p <= Pix_171;
    10'd4:  neuron_2_mul_6_p <= Pix_172;
    10'd5:  neuron_2_mul_6_p <= Pix_173;
    10'd6:  neuron_2_mul_6_p <= Pix_174;
    10'd7:  neuron_2_mul_6_p <= Pix_175;
    10'd8:  neuron_2_mul_6_p <= Pix_176;
    10'd9:  neuron_2_mul_6_p <= Pix_177;
    10'd10:  neuron_2_mul_6_p <= Pix_178;
    10'd11:  neuron_2_mul_6_p <= Pix_179;
    10'd12:  neuron_2_mul_6_p <= Pix_180;
    10'd13:  neuron_2_mul_6_p <= Pix_181;
    10'd14:  neuron_2_mul_6_p <= Pix_182;
    10'd15:  neuron_2_mul_6_p <= Pix_183;
    10'd16:  neuron_2_mul_6_p <= Pix_184;
    10'd17:  neuron_2_mul_6_p <= Pix_185;
    10'd18:  neuron_2_mul_6_p <= Pix_186;
    10'd19:  neuron_2_mul_6_p <= Pix_187;
    10'd20:  neuron_2_mul_6_p <= Pix_188;
    10'd21:  neuron_2_mul_6_p <= Pix_189;
    10'd22:  neuron_2_mul_6_p <= Pix_190;
    10'd23:  neuron_2_mul_6_p <= Pix_191;
    10'd24:  neuron_2_mul_6_p <= Pix_192;
    10'd25:  neuron_2_mul_6_p <= Pix_193;
    10'd26:  neuron_2_mul_6_p <= Pix_194;
    10'd27:  neuron_2_mul_6_p <= Pix_195;
    default: neuron_2_mul_6_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_7_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_7_p <= Pix_196;
    10'd1:  neuron_2_mul_7_p <= Pix_197;
    10'd2:  neuron_2_mul_7_p <= Pix_198;
    10'd3:  neuron_2_mul_7_p <= Pix_199;
    10'd4:  neuron_2_mul_7_p <= Pix_200;
    10'd5:  neuron_2_mul_7_p <= Pix_201;
    10'd6:  neuron_2_mul_7_p <= Pix_202;
    10'd7:  neuron_2_mul_7_p <= Pix_203;
    10'd8:  neuron_2_mul_7_p <= Pix_204;
    10'd9:  neuron_2_mul_7_p <= Pix_205;
    10'd10:  neuron_2_mul_7_p <= Pix_206;
    10'd11:  neuron_2_mul_7_p <= Pix_207;
    10'd12:  neuron_2_mul_7_p <= Pix_208;
    10'd13:  neuron_2_mul_7_p <= Pix_209;
    10'd14:  neuron_2_mul_7_p <= Pix_210;
    10'd15:  neuron_2_mul_7_p <= Pix_211;
    10'd16:  neuron_2_mul_7_p <= Pix_212;
    10'd17:  neuron_2_mul_7_p <= Pix_213;
    10'd18:  neuron_2_mul_7_p <= Pix_214;
    10'd19:  neuron_2_mul_7_p <= Pix_215;
    10'd20:  neuron_2_mul_7_p <= Pix_216;
    10'd21:  neuron_2_mul_7_p <= Pix_217;
    10'd22:  neuron_2_mul_7_p <= Pix_218;
    10'd23:  neuron_2_mul_7_p <= Pix_219;
    10'd24:  neuron_2_mul_7_p <= Pix_220;
    10'd25:  neuron_2_mul_7_p <= Pix_221;
    10'd26:  neuron_2_mul_7_p <= Pix_222;
    10'd27:  neuron_2_mul_7_p <= Pix_223;
    default: neuron_2_mul_7_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_8_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_8_p <= Pix_224;
    10'd1:  neuron_2_mul_8_p <= Pix_225;
    10'd2:  neuron_2_mul_8_p <= Pix_226;
    10'd3:  neuron_2_mul_8_p <= Pix_227;
    10'd4:  neuron_2_mul_8_p <= Pix_228;
    10'd5:  neuron_2_mul_8_p <= Pix_229;
    10'd6:  neuron_2_mul_8_p <= Pix_230;
    10'd7:  neuron_2_mul_8_p <= Pix_231;
    10'd8:  neuron_2_mul_8_p <= Pix_232;
    10'd9:  neuron_2_mul_8_p <= Pix_233;
    10'd10:  neuron_2_mul_8_p <= Pix_234;
    10'd11:  neuron_2_mul_8_p <= Pix_235;
    10'd12:  neuron_2_mul_8_p <= Pix_236;
    10'd13:  neuron_2_mul_8_p <= Pix_237;
    10'd14:  neuron_2_mul_8_p <= Pix_238;
    10'd15:  neuron_2_mul_8_p <= Pix_239;
    10'd16:  neuron_2_mul_8_p <= Pix_240;
    10'd17:  neuron_2_mul_8_p <= Pix_241;
    10'd18:  neuron_2_mul_8_p <= Pix_242;
    10'd19:  neuron_2_mul_8_p <= Pix_243;
    10'd20:  neuron_2_mul_8_p <= Pix_244;
    10'd21:  neuron_2_mul_8_p <= Pix_245;
    10'd22:  neuron_2_mul_8_p <= Pix_246;
    10'd23:  neuron_2_mul_8_p <= Pix_247;
    10'd24:  neuron_2_mul_8_p <= Pix_248;
    10'd25:  neuron_2_mul_8_p <= Pix_249;
    10'd26:  neuron_2_mul_8_p <= Pix_250;
    10'd27:  neuron_2_mul_8_p <= Pix_251;
    default: neuron_2_mul_8_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_9_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_9_p <= Pix_252;
    10'd1:  neuron_2_mul_9_p <= Pix_253;
    10'd2:  neuron_2_mul_9_p <= Pix_254;
    10'd3:  neuron_2_mul_9_p <= Pix_255;
    10'd4:  neuron_2_mul_9_p <= Pix_256;
    10'd5:  neuron_2_mul_9_p <= Pix_257;
    10'd6:  neuron_2_mul_9_p <= Pix_258;
    10'd7:  neuron_2_mul_9_p <= Pix_259;
    10'd8:  neuron_2_mul_9_p <= Pix_260;
    10'd9:  neuron_2_mul_9_p <= Pix_261;
    10'd10:  neuron_2_mul_9_p <= Pix_262;
    10'd11:  neuron_2_mul_9_p <= Pix_263;
    10'd12:  neuron_2_mul_9_p <= Pix_264;
    10'd13:  neuron_2_mul_9_p <= Pix_265;
    10'd14:  neuron_2_mul_9_p <= Pix_266;
    10'd15:  neuron_2_mul_9_p <= Pix_267;
    10'd16:  neuron_2_mul_9_p <= Pix_268;
    10'd17:  neuron_2_mul_9_p <= Pix_269;
    10'd18:  neuron_2_mul_9_p <= Pix_270;
    10'd19:  neuron_2_mul_9_p <= Pix_271;
    10'd20:  neuron_2_mul_9_p <= Pix_272;
    10'd21:  neuron_2_mul_9_p <= Pix_273;
    10'd22:  neuron_2_mul_9_p <= Pix_274;
    10'd23:  neuron_2_mul_9_p <= Pix_275;
    10'd24:  neuron_2_mul_9_p <= Pix_276;
    10'd25:  neuron_2_mul_9_p <= Pix_277;
    10'd26:  neuron_2_mul_9_p <= Pix_278;
    10'd27:  neuron_2_mul_9_p <= Pix_279;
    default: neuron_2_mul_9_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_10_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_10_p <= Pix_280;
    10'd1:  neuron_2_mul_10_p <= Pix_281;
    10'd2:  neuron_2_mul_10_p <= Pix_282;
    10'd3:  neuron_2_mul_10_p <= Pix_283;
    10'd4:  neuron_2_mul_10_p <= Pix_284;
    10'd5:  neuron_2_mul_10_p <= Pix_285;
    10'd6:  neuron_2_mul_10_p <= Pix_286;
    10'd7:  neuron_2_mul_10_p <= Pix_287;
    10'd8:  neuron_2_mul_10_p <= Pix_288;
    10'd9:  neuron_2_mul_10_p <= Pix_289;
    10'd10:  neuron_2_mul_10_p <= Pix_290;
    10'd11:  neuron_2_mul_10_p <= Pix_291;
    10'd12:  neuron_2_mul_10_p <= Pix_292;
    10'd13:  neuron_2_mul_10_p <= Pix_293;
    10'd14:  neuron_2_mul_10_p <= Pix_294;
    10'd15:  neuron_2_mul_10_p <= Pix_295;
    10'd16:  neuron_2_mul_10_p <= Pix_296;
    10'd17:  neuron_2_mul_10_p <= Pix_297;
    10'd18:  neuron_2_mul_10_p <= Pix_298;
    10'd19:  neuron_2_mul_10_p <= Pix_299;
    10'd20:  neuron_2_mul_10_p <= Pix_300;
    10'd21:  neuron_2_mul_10_p <= Pix_301;
    10'd22:  neuron_2_mul_10_p <= Pix_302;
    10'd23:  neuron_2_mul_10_p <= Pix_303;
    10'd24:  neuron_2_mul_10_p <= Pix_304;
    10'd25:  neuron_2_mul_10_p <= Pix_305;
    10'd26:  neuron_2_mul_10_p <= Pix_306;
    10'd27:  neuron_2_mul_10_p <= Pix_307;
    default: neuron_2_mul_10_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_11_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_11_p <= Pix_308;
    10'd1:  neuron_2_mul_11_p <= Pix_309;
    10'd2:  neuron_2_mul_11_p <= Pix_310;
    10'd3:  neuron_2_mul_11_p <= Pix_311;
    10'd4:  neuron_2_mul_11_p <= Pix_312;
    10'd5:  neuron_2_mul_11_p <= Pix_313;
    10'd6:  neuron_2_mul_11_p <= Pix_314;
    10'd7:  neuron_2_mul_11_p <= Pix_315;
    10'd8:  neuron_2_mul_11_p <= Pix_316;
    10'd9:  neuron_2_mul_11_p <= Pix_317;
    10'd10:  neuron_2_mul_11_p <= Pix_318;
    10'd11:  neuron_2_mul_11_p <= Pix_319;
    10'd12:  neuron_2_mul_11_p <= Pix_320;
    10'd13:  neuron_2_mul_11_p <= Pix_321;
    10'd14:  neuron_2_mul_11_p <= Pix_322;
    10'd15:  neuron_2_mul_11_p <= Pix_323;
    10'd16:  neuron_2_mul_11_p <= Pix_324;
    10'd17:  neuron_2_mul_11_p <= Pix_325;
    10'd18:  neuron_2_mul_11_p <= Pix_326;
    10'd19:  neuron_2_mul_11_p <= Pix_327;
    10'd20:  neuron_2_mul_11_p <= Pix_328;
    10'd21:  neuron_2_mul_11_p <= Pix_329;
    10'd22:  neuron_2_mul_11_p <= Pix_330;
    10'd23:  neuron_2_mul_11_p <= Pix_331;
    10'd24:  neuron_2_mul_11_p <= Pix_332;
    10'd25:  neuron_2_mul_11_p <= Pix_333;
    10'd26:  neuron_2_mul_11_p <= Pix_334;
    10'd27:  neuron_2_mul_11_p <= Pix_335;
    default: neuron_2_mul_11_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_12_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_12_p <= Pix_336;
    10'd1:  neuron_2_mul_12_p <= Pix_337;
    10'd2:  neuron_2_mul_12_p <= Pix_338;
    10'd3:  neuron_2_mul_12_p <= Pix_339;
    10'd4:  neuron_2_mul_12_p <= Pix_340;
    10'd5:  neuron_2_mul_12_p <= Pix_341;
    10'd6:  neuron_2_mul_12_p <= Pix_342;
    10'd7:  neuron_2_mul_12_p <= Pix_343;
    10'd8:  neuron_2_mul_12_p <= Pix_344;
    10'd9:  neuron_2_mul_12_p <= Pix_345;
    10'd10:  neuron_2_mul_12_p <= Pix_346;
    10'd11:  neuron_2_mul_12_p <= Pix_347;
    10'd12:  neuron_2_mul_12_p <= Pix_348;
    10'd13:  neuron_2_mul_12_p <= Pix_349;
    10'd14:  neuron_2_mul_12_p <= Pix_350;
    10'd15:  neuron_2_mul_12_p <= Pix_351;
    10'd16:  neuron_2_mul_12_p <= Pix_352;
    10'd17:  neuron_2_mul_12_p <= Pix_353;
    10'd18:  neuron_2_mul_12_p <= Pix_354;
    10'd19:  neuron_2_mul_12_p <= Pix_355;
    10'd20:  neuron_2_mul_12_p <= Pix_356;
    10'd21:  neuron_2_mul_12_p <= Pix_357;
    10'd22:  neuron_2_mul_12_p <= Pix_358;
    10'd23:  neuron_2_mul_12_p <= Pix_359;
    10'd24:  neuron_2_mul_12_p <= Pix_360;
    10'd25:  neuron_2_mul_12_p <= Pix_361;
    10'd26:  neuron_2_mul_12_p <= Pix_362;
    10'd27:  neuron_2_mul_12_p <= Pix_363;
    default: neuron_2_mul_12_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_13_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_13_p <= Pix_364;
    10'd1:  neuron_2_mul_13_p <= Pix_365;
    10'd2:  neuron_2_mul_13_p <= Pix_366;
    10'd3:  neuron_2_mul_13_p <= Pix_367;
    10'd4:  neuron_2_mul_13_p <= Pix_368;
    10'd5:  neuron_2_mul_13_p <= Pix_369;
    10'd6:  neuron_2_mul_13_p <= Pix_370;
    10'd7:  neuron_2_mul_13_p <= Pix_371;
    10'd8:  neuron_2_mul_13_p <= Pix_372;
    10'd9:  neuron_2_mul_13_p <= Pix_373;
    10'd10:  neuron_2_mul_13_p <= Pix_374;
    10'd11:  neuron_2_mul_13_p <= Pix_375;
    10'd12:  neuron_2_mul_13_p <= Pix_376;
    10'd13:  neuron_2_mul_13_p <= Pix_377;
    10'd14:  neuron_2_mul_13_p <= Pix_378;
    10'd15:  neuron_2_mul_13_p <= Pix_379;
    10'd16:  neuron_2_mul_13_p <= Pix_380;
    10'd17:  neuron_2_mul_13_p <= Pix_381;
    10'd18:  neuron_2_mul_13_p <= Pix_382;
    10'd19:  neuron_2_mul_13_p <= Pix_383;
    10'd20:  neuron_2_mul_13_p <= Pix_384;
    10'd21:  neuron_2_mul_13_p <= Pix_385;
    10'd22:  neuron_2_mul_13_p <= Pix_386;
    10'd23:  neuron_2_mul_13_p <= Pix_387;
    10'd24:  neuron_2_mul_13_p <= Pix_388;
    10'd25:  neuron_2_mul_13_p <= Pix_389;
    10'd26:  neuron_2_mul_13_p <= Pix_390;
    10'd27:  neuron_2_mul_13_p <= Pix_391;
    default: neuron_2_mul_13_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_14_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_14_p <= Pix_392;
    10'd1:  neuron_2_mul_14_p <= Pix_393;
    10'd2:  neuron_2_mul_14_p <= Pix_394;
    10'd3:  neuron_2_mul_14_p <= Pix_395;
    10'd4:  neuron_2_mul_14_p <= Pix_396;
    10'd5:  neuron_2_mul_14_p <= Pix_397;
    10'd6:  neuron_2_mul_14_p <= Pix_398;
    10'd7:  neuron_2_mul_14_p <= Pix_399;
    10'd8:  neuron_2_mul_14_p <= Pix_400;
    10'd9:  neuron_2_mul_14_p <= Pix_401;
    10'd10:  neuron_2_mul_14_p <= Pix_402;
    10'd11:  neuron_2_mul_14_p <= Pix_403;
    10'd12:  neuron_2_mul_14_p <= Pix_404;
    10'd13:  neuron_2_mul_14_p <= Pix_405;
    10'd14:  neuron_2_mul_14_p <= Pix_406;
    10'd15:  neuron_2_mul_14_p <= Pix_407;
    10'd16:  neuron_2_mul_14_p <= Pix_408;
    10'd17:  neuron_2_mul_14_p <= Pix_409;
    10'd18:  neuron_2_mul_14_p <= Pix_410;
    10'd19:  neuron_2_mul_14_p <= Pix_411;
    10'd20:  neuron_2_mul_14_p <= Pix_412;
    10'd21:  neuron_2_mul_14_p <= Pix_413;
    10'd22:  neuron_2_mul_14_p <= Pix_414;
    10'd23:  neuron_2_mul_14_p <= Pix_415;
    10'd24:  neuron_2_mul_14_p <= Pix_416;
    10'd25:  neuron_2_mul_14_p <= Pix_417;
    10'd26:  neuron_2_mul_14_p <= Pix_418;
    10'd27:  neuron_2_mul_14_p <= Pix_419;
    default: neuron_2_mul_14_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_15_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_15_p <= Pix_420;
    10'd1:  neuron_2_mul_15_p <= Pix_421;
    10'd2:  neuron_2_mul_15_p <= Pix_422;
    10'd3:  neuron_2_mul_15_p <= Pix_423;
    10'd4:  neuron_2_mul_15_p <= Pix_424;
    10'd5:  neuron_2_mul_15_p <= Pix_425;
    10'd6:  neuron_2_mul_15_p <= Pix_426;
    10'd7:  neuron_2_mul_15_p <= Pix_427;
    10'd8:  neuron_2_mul_15_p <= Pix_428;
    10'd9:  neuron_2_mul_15_p <= Pix_429;
    10'd10:  neuron_2_mul_15_p <= Pix_430;
    10'd11:  neuron_2_mul_15_p <= Pix_431;
    10'd12:  neuron_2_mul_15_p <= Pix_432;
    10'd13:  neuron_2_mul_15_p <= Pix_433;
    10'd14:  neuron_2_mul_15_p <= Pix_434;
    10'd15:  neuron_2_mul_15_p <= Pix_435;
    10'd16:  neuron_2_mul_15_p <= Pix_436;
    10'd17:  neuron_2_mul_15_p <= Pix_437;
    10'd18:  neuron_2_mul_15_p <= Pix_438;
    10'd19:  neuron_2_mul_15_p <= Pix_439;
    10'd20:  neuron_2_mul_15_p <= Pix_440;
    10'd21:  neuron_2_mul_15_p <= Pix_441;
    10'd22:  neuron_2_mul_15_p <= Pix_442;
    10'd23:  neuron_2_mul_15_p <= Pix_443;
    10'd24:  neuron_2_mul_15_p <= Pix_444;
    10'd25:  neuron_2_mul_15_p <= Pix_445;
    10'd26:  neuron_2_mul_15_p <= Pix_446;
    10'd27:  neuron_2_mul_15_p <= Pix_447;
    default: neuron_2_mul_15_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_16_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_16_p <= Pix_448;
    10'd1:  neuron_2_mul_16_p <= Pix_449;
    10'd2:  neuron_2_mul_16_p <= Pix_450;
    10'd3:  neuron_2_mul_16_p <= Pix_451;
    10'd4:  neuron_2_mul_16_p <= Pix_452;
    10'd5:  neuron_2_mul_16_p <= Pix_453;
    10'd6:  neuron_2_mul_16_p <= Pix_454;
    10'd7:  neuron_2_mul_16_p <= Pix_455;
    10'd8:  neuron_2_mul_16_p <= Pix_456;
    10'd9:  neuron_2_mul_16_p <= Pix_457;
    10'd10:  neuron_2_mul_16_p <= Pix_458;
    10'd11:  neuron_2_mul_16_p <= Pix_459;
    10'd12:  neuron_2_mul_16_p <= Pix_460;
    10'd13:  neuron_2_mul_16_p <= Pix_461;
    10'd14:  neuron_2_mul_16_p <= Pix_462;
    10'd15:  neuron_2_mul_16_p <= Pix_463;
    10'd16:  neuron_2_mul_16_p <= Pix_464;
    10'd17:  neuron_2_mul_16_p <= Pix_465;
    10'd18:  neuron_2_mul_16_p <= Pix_466;
    10'd19:  neuron_2_mul_16_p <= Pix_467;
    10'd20:  neuron_2_mul_16_p <= Pix_468;
    10'd21:  neuron_2_mul_16_p <= Pix_469;
    10'd22:  neuron_2_mul_16_p <= Pix_470;
    10'd23:  neuron_2_mul_16_p <= Pix_471;
    10'd24:  neuron_2_mul_16_p <= Pix_472;
    10'd25:  neuron_2_mul_16_p <= Pix_473;
    10'd26:  neuron_2_mul_16_p <= Pix_474;
    10'd27:  neuron_2_mul_16_p <= Pix_475;
    default: neuron_2_mul_16_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_17_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_17_p <= Pix_476;
    10'd1:  neuron_2_mul_17_p <= Pix_477;
    10'd2:  neuron_2_mul_17_p <= Pix_478;
    10'd3:  neuron_2_mul_17_p <= Pix_479;
    10'd4:  neuron_2_mul_17_p <= Pix_480;
    10'd5:  neuron_2_mul_17_p <= Pix_481;
    10'd6:  neuron_2_mul_17_p <= Pix_482;
    10'd7:  neuron_2_mul_17_p <= Pix_483;
    10'd8:  neuron_2_mul_17_p <= Pix_484;
    10'd9:  neuron_2_mul_17_p <= Pix_485;
    10'd10:  neuron_2_mul_17_p <= Pix_486;
    10'd11:  neuron_2_mul_17_p <= Pix_487;
    10'd12:  neuron_2_mul_17_p <= Pix_488;
    10'd13:  neuron_2_mul_17_p <= Pix_489;
    10'd14:  neuron_2_mul_17_p <= Pix_490;
    10'd15:  neuron_2_mul_17_p <= Pix_491;
    10'd16:  neuron_2_mul_17_p <= Pix_492;
    10'd17:  neuron_2_mul_17_p <= Pix_493;
    10'd18:  neuron_2_mul_17_p <= Pix_494;
    10'd19:  neuron_2_mul_17_p <= Pix_495;
    10'd20:  neuron_2_mul_17_p <= Pix_496;
    10'd21:  neuron_2_mul_17_p <= Pix_497;
    10'd22:  neuron_2_mul_17_p <= Pix_498;
    10'd23:  neuron_2_mul_17_p <= Pix_499;
    10'd24:  neuron_2_mul_17_p <= Pix_500;
    10'd25:  neuron_2_mul_17_p <= Pix_501;
    10'd26:  neuron_2_mul_17_p <= Pix_502;
    10'd27:  neuron_2_mul_17_p <= Pix_503;
    default: neuron_2_mul_17_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_18_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_18_p <= Pix_504;
    10'd1:  neuron_2_mul_18_p <= Pix_505;
    10'd2:  neuron_2_mul_18_p <= Pix_506;
    10'd3:  neuron_2_mul_18_p <= Pix_507;
    10'd4:  neuron_2_mul_18_p <= Pix_508;
    10'd5:  neuron_2_mul_18_p <= Pix_509;
    10'd6:  neuron_2_mul_18_p <= Pix_510;
    10'd7:  neuron_2_mul_18_p <= Pix_511;
    10'd8:  neuron_2_mul_18_p <= Pix_512;
    10'd9:  neuron_2_mul_18_p <= Pix_513;
    10'd10:  neuron_2_mul_18_p <= Pix_514;
    10'd11:  neuron_2_mul_18_p <= Pix_515;
    10'd12:  neuron_2_mul_18_p <= Pix_516;
    10'd13:  neuron_2_mul_18_p <= Pix_517;
    10'd14:  neuron_2_mul_18_p <= Pix_518;
    10'd15:  neuron_2_mul_18_p <= Pix_519;
    10'd16:  neuron_2_mul_18_p <= Pix_520;
    10'd17:  neuron_2_mul_18_p <= Pix_521;
    10'd18:  neuron_2_mul_18_p <= Pix_522;
    10'd19:  neuron_2_mul_18_p <= Pix_523;
    10'd20:  neuron_2_mul_18_p <= Pix_524;
    10'd21:  neuron_2_mul_18_p <= Pix_525;
    10'd22:  neuron_2_mul_18_p <= Pix_526;
    10'd23:  neuron_2_mul_18_p <= Pix_527;
    10'd24:  neuron_2_mul_18_p <= Pix_528;
    10'd25:  neuron_2_mul_18_p <= Pix_529;
    10'd26:  neuron_2_mul_18_p <= Pix_530;
    10'd27:  neuron_2_mul_18_p <= Pix_531;
    default: neuron_2_mul_18_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_19_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_19_p <= Pix_532;
    10'd1:  neuron_2_mul_19_p <= Pix_533;
    10'd2:  neuron_2_mul_19_p <= Pix_534;
    10'd3:  neuron_2_mul_19_p <= Pix_535;
    10'd4:  neuron_2_mul_19_p <= Pix_536;
    10'd5:  neuron_2_mul_19_p <= Pix_537;
    10'd6:  neuron_2_mul_19_p <= Pix_538;
    10'd7:  neuron_2_mul_19_p <= Pix_539;
    10'd8:  neuron_2_mul_19_p <= Pix_540;
    10'd9:  neuron_2_mul_19_p <= Pix_541;
    10'd10:  neuron_2_mul_19_p <= Pix_542;
    10'd11:  neuron_2_mul_19_p <= Pix_543;
    10'd12:  neuron_2_mul_19_p <= Pix_544;
    10'd13:  neuron_2_mul_19_p <= Pix_545;
    10'd14:  neuron_2_mul_19_p <= Pix_546;
    10'd15:  neuron_2_mul_19_p <= Pix_547;
    10'd16:  neuron_2_mul_19_p <= Pix_548;
    10'd17:  neuron_2_mul_19_p <= Pix_549;
    10'd18:  neuron_2_mul_19_p <= Pix_550;
    10'd19:  neuron_2_mul_19_p <= Pix_551;
    10'd20:  neuron_2_mul_19_p <= Pix_552;
    10'd21:  neuron_2_mul_19_p <= Pix_553;
    10'd22:  neuron_2_mul_19_p <= Pix_554;
    10'd23:  neuron_2_mul_19_p <= Pix_555;
    10'd24:  neuron_2_mul_19_p <= Pix_556;
    10'd25:  neuron_2_mul_19_p <= Pix_557;
    10'd26:  neuron_2_mul_19_p <= Pix_558;
    10'd27:  neuron_2_mul_19_p <= Pix_559;
    default: neuron_2_mul_19_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_20_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_20_p <= Pix_560;
    10'd1:  neuron_2_mul_20_p <= Pix_561;
    10'd2:  neuron_2_mul_20_p <= Pix_562;
    10'd3:  neuron_2_mul_20_p <= Pix_563;
    10'd4:  neuron_2_mul_20_p <= Pix_564;
    10'd5:  neuron_2_mul_20_p <= Pix_565;
    10'd6:  neuron_2_mul_20_p <= Pix_566;
    10'd7:  neuron_2_mul_20_p <= Pix_567;
    10'd8:  neuron_2_mul_20_p <= Pix_568;
    10'd9:  neuron_2_mul_20_p <= Pix_569;
    10'd10:  neuron_2_mul_20_p <= Pix_570;
    10'd11:  neuron_2_mul_20_p <= Pix_571;
    10'd12:  neuron_2_mul_20_p <= Pix_572;
    10'd13:  neuron_2_mul_20_p <= Pix_573;
    10'd14:  neuron_2_mul_20_p <= Pix_574;
    10'd15:  neuron_2_mul_20_p <= Pix_575;
    10'd16:  neuron_2_mul_20_p <= Pix_576;
    10'd17:  neuron_2_mul_20_p <= Pix_577;
    10'd18:  neuron_2_mul_20_p <= Pix_578;
    10'd19:  neuron_2_mul_20_p <= Pix_579;
    10'd20:  neuron_2_mul_20_p <= Pix_580;
    10'd21:  neuron_2_mul_20_p <= Pix_581;
    10'd22:  neuron_2_mul_20_p <= Pix_582;
    10'd23:  neuron_2_mul_20_p <= Pix_583;
    10'd24:  neuron_2_mul_20_p <= Pix_584;
    10'd25:  neuron_2_mul_20_p <= Pix_585;
    10'd26:  neuron_2_mul_20_p <= Pix_586;
    10'd27:  neuron_2_mul_20_p <= Pix_587;
    default: neuron_2_mul_20_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_21_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_21_p <= Pix_588;
    10'd1:  neuron_2_mul_21_p <= Pix_589;
    10'd2:  neuron_2_mul_21_p <= Pix_590;
    10'd3:  neuron_2_mul_21_p <= Pix_591;
    10'd4:  neuron_2_mul_21_p <= Pix_592;
    10'd5:  neuron_2_mul_21_p <= Pix_593;
    10'd6:  neuron_2_mul_21_p <= Pix_594;
    10'd7:  neuron_2_mul_21_p <= Pix_595;
    10'd8:  neuron_2_mul_21_p <= Pix_596;
    10'd9:  neuron_2_mul_21_p <= Pix_597;
    10'd10:  neuron_2_mul_21_p <= Pix_598;
    10'd11:  neuron_2_mul_21_p <= Pix_599;
    10'd12:  neuron_2_mul_21_p <= Pix_600;
    10'd13:  neuron_2_mul_21_p <= Pix_601;
    10'd14:  neuron_2_mul_21_p <= Pix_602;
    10'd15:  neuron_2_mul_21_p <= Pix_603;
    10'd16:  neuron_2_mul_21_p <= Pix_604;
    10'd17:  neuron_2_mul_21_p <= Pix_605;
    10'd18:  neuron_2_mul_21_p <= Pix_606;
    10'd19:  neuron_2_mul_21_p <= Pix_607;
    10'd20:  neuron_2_mul_21_p <= Pix_608;
    10'd21:  neuron_2_mul_21_p <= Pix_609;
    10'd22:  neuron_2_mul_21_p <= Pix_610;
    10'd23:  neuron_2_mul_21_p <= Pix_611;
    10'd24:  neuron_2_mul_21_p <= Pix_612;
    10'd25:  neuron_2_mul_21_p <= Pix_613;
    10'd26:  neuron_2_mul_21_p <= Pix_614;
    10'd27:  neuron_2_mul_21_p <= Pix_615;
    default: neuron_2_mul_21_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_22_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_22_p <= Pix_616;
    10'd1:  neuron_2_mul_22_p <= Pix_617;
    10'd2:  neuron_2_mul_22_p <= Pix_618;
    10'd3:  neuron_2_mul_22_p <= Pix_619;
    10'd4:  neuron_2_mul_22_p <= Pix_620;
    10'd5:  neuron_2_mul_22_p <= Pix_621;
    10'd6:  neuron_2_mul_22_p <= Pix_622;
    10'd7:  neuron_2_mul_22_p <= Pix_623;
    10'd8:  neuron_2_mul_22_p <= Pix_624;
    10'd9:  neuron_2_mul_22_p <= Pix_625;
    10'd10:  neuron_2_mul_22_p <= Pix_626;
    10'd11:  neuron_2_mul_22_p <= Pix_627;
    10'd12:  neuron_2_mul_22_p <= Pix_628;
    10'd13:  neuron_2_mul_22_p <= Pix_629;
    10'd14:  neuron_2_mul_22_p <= Pix_630;
    10'd15:  neuron_2_mul_22_p <= Pix_631;
    10'd16:  neuron_2_mul_22_p <= Pix_632;
    10'd17:  neuron_2_mul_22_p <= Pix_633;
    10'd18:  neuron_2_mul_22_p <= Pix_634;
    10'd19:  neuron_2_mul_22_p <= Pix_635;
    10'd20:  neuron_2_mul_22_p <= Pix_636;
    10'd21:  neuron_2_mul_22_p <= Pix_637;
    10'd22:  neuron_2_mul_22_p <= Pix_638;
    10'd23:  neuron_2_mul_22_p <= Pix_639;
    10'd24:  neuron_2_mul_22_p <= Pix_640;
    10'd25:  neuron_2_mul_22_p <= Pix_641;
    10'd26:  neuron_2_mul_22_p <= Pix_642;
    10'd27:  neuron_2_mul_22_p <= Pix_643;
    default: neuron_2_mul_22_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_23_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_23_p <= Pix_644;
    10'd1:  neuron_2_mul_23_p <= Pix_645;
    10'd2:  neuron_2_mul_23_p <= Pix_646;
    10'd3:  neuron_2_mul_23_p <= Pix_647;
    10'd4:  neuron_2_mul_23_p <= Pix_648;
    10'd5:  neuron_2_mul_23_p <= Pix_649;
    10'd6:  neuron_2_mul_23_p <= Pix_650;
    10'd7:  neuron_2_mul_23_p <= Pix_651;
    10'd8:  neuron_2_mul_23_p <= Pix_652;
    10'd9:  neuron_2_mul_23_p <= Pix_653;
    10'd10:  neuron_2_mul_23_p <= Pix_654;
    10'd11:  neuron_2_mul_23_p <= Pix_655;
    10'd12:  neuron_2_mul_23_p <= Pix_656;
    10'd13:  neuron_2_mul_23_p <= Pix_657;
    10'd14:  neuron_2_mul_23_p <= Pix_658;
    10'd15:  neuron_2_mul_23_p <= Pix_659;
    10'd16:  neuron_2_mul_23_p <= Pix_660;
    10'd17:  neuron_2_mul_23_p <= Pix_661;
    10'd18:  neuron_2_mul_23_p <= Pix_662;
    10'd19:  neuron_2_mul_23_p <= Pix_663;
    10'd20:  neuron_2_mul_23_p <= Pix_664;
    10'd21:  neuron_2_mul_23_p <= Pix_665;
    10'd22:  neuron_2_mul_23_p <= Pix_666;
    10'd23:  neuron_2_mul_23_p <= Pix_667;
    10'd24:  neuron_2_mul_23_p <= Pix_668;
    10'd25:  neuron_2_mul_23_p <= Pix_669;
    10'd26:  neuron_2_mul_23_p <= Pix_670;
    10'd27:  neuron_2_mul_23_p <= Pix_671;
    default: neuron_2_mul_23_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_24_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_24_p <= Pix_672;
    10'd1:  neuron_2_mul_24_p <= Pix_673;
    10'd2:  neuron_2_mul_24_p <= Pix_674;
    10'd3:  neuron_2_mul_24_p <= Pix_675;
    10'd4:  neuron_2_mul_24_p <= Pix_676;
    10'd5:  neuron_2_mul_24_p <= Pix_677;
    10'd6:  neuron_2_mul_24_p <= Pix_678;
    10'd7:  neuron_2_mul_24_p <= Pix_679;
    10'd8:  neuron_2_mul_24_p <= Pix_680;
    10'd9:  neuron_2_mul_24_p <= Pix_681;
    10'd10:  neuron_2_mul_24_p <= Pix_682;
    10'd11:  neuron_2_mul_24_p <= Pix_683;
    10'd12:  neuron_2_mul_24_p <= Pix_684;
    10'd13:  neuron_2_mul_24_p <= Pix_685;
    10'd14:  neuron_2_mul_24_p <= Pix_686;
    10'd15:  neuron_2_mul_24_p <= Pix_687;
    10'd16:  neuron_2_mul_24_p <= Pix_688;
    10'd17:  neuron_2_mul_24_p <= Pix_689;
    10'd18:  neuron_2_mul_24_p <= Pix_690;
    10'd19:  neuron_2_mul_24_p <= Pix_691;
    10'd20:  neuron_2_mul_24_p <= Pix_692;
    10'd21:  neuron_2_mul_24_p <= Pix_693;
    10'd22:  neuron_2_mul_24_p <= Pix_694;
    10'd23:  neuron_2_mul_24_p <= Pix_695;
    10'd24:  neuron_2_mul_24_p <= Pix_696;
    10'd25:  neuron_2_mul_24_p <= Pix_697;
    10'd26:  neuron_2_mul_24_p <= Pix_698;
    10'd27:  neuron_2_mul_24_p <= Pix_699;
    default: neuron_2_mul_24_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_25_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_25_p <= Pix_700;
    10'd1:  neuron_2_mul_25_p <= Pix_701;
    10'd2:  neuron_2_mul_25_p <= Pix_702;
    10'd3:  neuron_2_mul_25_p <= Pix_703;
    10'd4:  neuron_2_mul_25_p <= Pix_704;
    10'd5:  neuron_2_mul_25_p <= Pix_705;
    10'd6:  neuron_2_mul_25_p <= Pix_706;
    10'd7:  neuron_2_mul_25_p <= Pix_707;
    10'd8:  neuron_2_mul_25_p <= Pix_708;
    10'd9:  neuron_2_mul_25_p <= Pix_709;
    10'd10:  neuron_2_mul_25_p <= Pix_710;
    10'd11:  neuron_2_mul_25_p <= Pix_711;
    10'd12:  neuron_2_mul_25_p <= Pix_712;
    10'd13:  neuron_2_mul_25_p <= Pix_713;
    10'd14:  neuron_2_mul_25_p <= Pix_714;
    10'd15:  neuron_2_mul_25_p <= Pix_715;
    10'd16:  neuron_2_mul_25_p <= Pix_716;
    10'd17:  neuron_2_mul_25_p <= Pix_717;
    10'd18:  neuron_2_mul_25_p <= Pix_718;
    10'd19:  neuron_2_mul_25_p <= Pix_719;
    10'd20:  neuron_2_mul_25_p <= Pix_720;
    10'd21:  neuron_2_mul_25_p <= Pix_721;
    10'd22:  neuron_2_mul_25_p <= Pix_722;
    10'd23:  neuron_2_mul_25_p <= Pix_723;
    10'd24:  neuron_2_mul_25_p <= Pix_724;
    10'd25:  neuron_2_mul_25_p <= Pix_725;
    10'd26:  neuron_2_mul_25_p <= Pix_726;
    10'd27:  neuron_2_mul_25_p <= Pix_727;
    default: neuron_2_mul_25_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_26_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_26_p <= Pix_728;
    10'd1:  neuron_2_mul_26_p <= Pix_729;
    10'd2:  neuron_2_mul_26_p <= Pix_730;
    10'd3:  neuron_2_mul_26_p <= Pix_731;
    10'd4:  neuron_2_mul_26_p <= Pix_732;
    10'd5:  neuron_2_mul_26_p <= Pix_733;
    10'd6:  neuron_2_mul_26_p <= Pix_734;
    10'd7:  neuron_2_mul_26_p <= Pix_735;
    10'd8:  neuron_2_mul_26_p <= Pix_736;
    10'd9:  neuron_2_mul_26_p <= Pix_737;
    10'd10:  neuron_2_mul_26_p <= Pix_738;
    10'd11:  neuron_2_mul_26_p <= Pix_739;
    10'd12:  neuron_2_mul_26_p <= Pix_740;
    10'd13:  neuron_2_mul_26_p <= Pix_741;
    10'd14:  neuron_2_mul_26_p <= Pix_742;
    10'd15:  neuron_2_mul_26_p <= Pix_743;
    10'd16:  neuron_2_mul_26_p <= Pix_744;
    10'd17:  neuron_2_mul_26_p <= Pix_745;
    10'd18:  neuron_2_mul_26_p <= Pix_746;
    10'd19:  neuron_2_mul_26_p <= Pix_747;
    10'd20:  neuron_2_mul_26_p <= Pix_748;
    10'd21:  neuron_2_mul_26_p <= Pix_749;
    10'd22:  neuron_2_mul_26_p <= Pix_750;
    10'd23:  neuron_2_mul_26_p <= Pix_751;
    10'd24:  neuron_2_mul_26_p <= Pix_752;
    10'd25:  neuron_2_mul_26_p <= Pix_753;
    10'd26:  neuron_2_mul_26_p <= Pix_754;
    10'd27:  neuron_2_mul_26_p <= Pix_755;
    default: neuron_2_mul_26_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_2_mul_27_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_2_mul_27_p <= Pix_756;
    10'd1:  neuron_2_mul_27_p <= Pix_757;
    10'd2:  neuron_2_mul_27_p <= Pix_758;
    10'd3:  neuron_2_mul_27_p <= Pix_759;
    10'd4:  neuron_2_mul_27_p <= Pix_760;
    10'd5:  neuron_2_mul_27_p <= Pix_761;
    10'd6:  neuron_2_mul_27_p <= Pix_762;
    10'd7:  neuron_2_mul_27_p <= Pix_763;
    10'd8:  neuron_2_mul_27_p <= Pix_764;
    10'd9:  neuron_2_mul_27_p <= Pix_765;
    10'd10:  neuron_2_mul_27_p <= Pix_766;
    10'd11:  neuron_2_mul_27_p <= Pix_767;
    10'd12:  neuron_2_mul_27_p <= Pix_768;
    10'd13:  neuron_2_mul_27_p <= Pix_769;
    10'd14:  neuron_2_mul_27_p <= Pix_770;
    10'd15:  neuron_2_mul_27_p <= Pix_771;
    10'd16:  neuron_2_mul_27_p <= Pix_772;
    10'd17:  neuron_2_mul_27_p <= Pix_773;
    10'd18:  neuron_2_mul_27_p <= Pix_774;
    10'd19:  neuron_2_mul_27_p <= Pix_775;
    10'd20:  neuron_2_mul_27_p <= Pix_776;
    10'd21:  neuron_2_mul_27_p <= Pix_777;
    10'd22:  neuron_2_mul_27_p <= Pix_778;
    10'd23:  neuron_2_mul_27_p <= Pix_779;
    10'd24:  neuron_2_mul_27_p <= Pix_780;
    10'd25:  neuron_2_mul_27_p <= Pix_781;
    10'd26:  neuron_2_mul_27_p <= Pix_782;
    10'd27:  neuron_2_mul_27_p <= Pix_783;
    default: neuron_2_mul_27_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_0_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_0_p <= Pix_0;
    10'd1:  neuron_3_mul_0_p <= Pix_1;
    10'd2:  neuron_3_mul_0_p <= Pix_2;
    10'd3:  neuron_3_mul_0_p <= Pix_3;
    10'd4:  neuron_3_mul_0_p <= Pix_4;
    10'd5:  neuron_3_mul_0_p <= Pix_5;
    10'd6:  neuron_3_mul_0_p <= Pix_6;
    10'd7:  neuron_3_mul_0_p <= Pix_7;
    10'd8:  neuron_3_mul_0_p <= Pix_8;
    10'd9:  neuron_3_mul_0_p <= Pix_9;
    10'd10:  neuron_3_mul_0_p <= Pix_10;
    10'd11:  neuron_3_mul_0_p <= Pix_11;
    10'd12:  neuron_3_mul_0_p <= Pix_12;
    10'd13:  neuron_3_mul_0_p <= Pix_13;
    10'd14:  neuron_3_mul_0_p <= Pix_14;
    10'd15:  neuron_3_mul_0_p <= Pix_15;
    10'd16:  neuron_3_mul_0_p <= Pix_16;
    10'd17:  neuron_3_mul_0_p <= Pix_17;
    10'd18:  neuron_3_mul_0_p <= Pix_18;
    10'd19:  neuron_3_mul_0_p <= Pix_19;
    10'd20:  neuron_3_mul_0_p <= Pix_20;
    10'd21:  neuron_3_mul_0_p <= Pix_21;
    10'd22:  neuron_3_mul_0_p <= Pix_22;
    10'd23:  neuron_3_mul_0_p <= Pix_23;
    10'd24:  neuron_3_mul_0_p <= Pix_24;
    10'd25:  neuron_3_mul_0_p <= Pix_25;
    10'd26:  neuron_3_mul_0_p <= Pix_26;
    10'd27:  neuron_3_mul_0_p <= Pix_27;
    default: neuron_3_mul_0_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_1_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_1_p <= Pix_28;
    10'd1:  neuron_3_mul_1_p <= Pix_29;
    10'd2:  neuron_3_mul_1_p <= Pix_30;
    10'd3:  neuron_3_mul_1_p <= Pix_31;
    10'd4:  neuron_3_mul_1_p <= Pix_32;
    10'd5:  neuron_3_mul_1_p <= Pix_33;
    10'd6:  neuron_3_mul_1_p <= Pix_34;
    10'd7:  neuron_3_mul_1_p <= Pix_35;
    10'd8:  neuron_3_mul_1_p <= Pix_36;
    10'd9:  neuron_3_mul_1_p <= Pix_37;
    10'd10:  neuron_3_mul_1_p <= Pix_38;
    10'd11:  neuron_3_mul_1_p <= Pix_39;
    10'd12:  neuron_3_mul_1_p <= Pix_40;
    10'd13:  neuron_3_mul_1_p <= Pix_41;
    10'd14:  neuron_3_mul_1_p <= Pix_42;
    10'd15:  neuron_3_mul_1_p <= Pix_43;
    10'd16:  neuron_3_mul_1_p <= Pix_44;
    10'd17:  neuron_3_mul_1_p <= Pix_45;
    10'd18:  neuron_3_mul_1_p <= Pix_46;
    10'd19:  neuron_3_mul_1_p <= Pix_47;
    10'd20:  neuron_3_mul_1_p <= Pix_48;
    10'd21:  neuron_3_mul_1_p <= Pix_49;
    10'd22:  neuron_3_mul_1_p <= Pix_50;
    10'd23:  neuron_3_mul_1_p <= Pix_51;
    10'd24:  neuron_3_mul_1_p <= Pix_52;
    10'd25:  neuron_3_mul_1_p <= Pix_53;
    10'd26:  neuron_3_mul_1_p <= Pix_54;
    10'd27:  neuron_3_mul_1_p <= Pix_55;
    default: neuron_3_mul_1_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_2_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_2_p <= Pix_56;
    10'd1:  neuron_3_mul_2_p <= Pix_57;
    10'd2:  neuron_3_mul_2_p <= Pix_58;
    10'd3:  neuron_3_mul_2_p <= Pix_59;
    10'd4:  neuron_3_mul_2_p <= Pix_60;
    10'd5:  neuron_3_mul_2_p <= Pix_61;
    10'd6:  neuron_3_mul_2_p <= Pix_62;
    10'd7:  neuron_3_mul_2_p <= Pix_63;
    10'd8:  neuron_3_mul_2_p <= Pix_64;
    10'd9:  neuron_3_mul_2_p <= Pix_65;
    10'd10:  neuron_3_mul_2_p <= Pix_66;
    10'd11:  neuron_3_mul_2_p <= Pix_67;
    10'd12:  neuron_3_mul_2_p <= Pix_68;
    10'd13:  neuron_3_mul_2_p <= Pix_69;
    10'd14:  neuron_3_mul_2_p <= Pix_70;
    10'd15:  neuron_3_mul_2_p <= Pix_71;
    10'd16:  neuron_3_mul_2_p <= Pix_72;
    10'd17:  neuron_3_mul_2_p <= Pix_73;
    10'd18:  neuron_3_mul_2_p <= Pix_74;
    10'd19:  neuron_3_mul_2_p <= Pix_75;
    10'd20:  neuron_3_mul_2_p <= Pix_76;
    10'd21:  neuron_3_mul_2_p <= Pix_77;
    10'd22:  neuron_3_mul_2_p <= Pix_78;
    10'd23:  neuron_3_mul_2_p <= Pix_79;
    10'd24:  neuron_3_mul_2_p <= Pix_80;
    10'd25:  neuron_3_mul_2_p <= Pix_81;
    10'd26:  neuron_3_mul_2_p <= Pix_82;
    10'd27:  neuron_3_mul_2_p <= Pix_83;
    default: neuron_3_mul_2_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_3_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_3_p <= Pix_84;
    10'd1:  neuron_3_mul_3_p <= Pix_85;
    10'd2:  neuron_3_mul_3_p <= Pix_86;
    10'd3:  neuron_3_mul_3_p <= Pix_87;
    10'd4:  neuron_3_mul_3_p <= Pix_88;
    10'd5:  neuron_3_mul_3_p <= Pix_89;
    10'd6:  neuron_3_mul_3_p <= Pix_90;
    10'd7:  neuron_3_mul_3_p <= Pix_91;
    10'd8:  neuron_3_mul_3_p <= Pix_92;
    10'd9:  neuron_3_mul_3_p <= Pix_93;
    10'd10:  neuron_3_mul_3_p <= Pix_94;
    10'd11:  neuron_3_mul_3_p <= Pix_95;
    10'd12:  neuron_3_mul_3_p <= Pix_96;
    10'd13:  neuron_3_mul_3_p <= Pix_97;
    10'd14:  neuron_3_mul_3_p <= Pix_98;
    10'd15:  neuron_3_mul_3_p <= Pix_99;
    10'd16:  neuron_3_mul_3_p <= Pix_100;
    10'd17:  neuron_3_mul_3_p <= Pix_101;
    10'd18:  neuron_3_mul_3_p <= Pix_102;
    10'd19:  neuron_3_mul_3_p <= Pix_103;
    10'd20:  neuron_3_mul_3_p <= Pix_104;
    10'd21:  neuron_3_mul_3_p <= Pix_105;
    10'd22:  neuron_3_mul_3_p <= Pix_106;
    10'd23:  neuron_3_mul_3_p <= Pix_107;
    10'd24:  neuron_3_mul_3_p <= Pix_108;
    10'd25:  neuron_3_mul_3_p <= Pix_109;
    10'd26:  neuron_3_mul_3_p <= Pix_110;
    10'd27:  neuron_3_mul_3_p <= Pix_111;
    default: neuron_3_mul_3_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_4_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_4_p <= Pix_112;
    10'd1:  neuron_3_mul_4_p <= Pix_113;
    10'd2:  neuron_3_mul_4_p <= Pix_114;
    10'd3:  neuron_3_mul_4_p <= Pix_115;
    10'd4:  neuron_3_mul_4_p <= Pix_116;
    10'd5:  neuron_3_mul_4_p <= Pix_117;
    10'd6:  neuron_3_mul_4_p <= Pix_118;
    10'd7:  neuron_3_mul_4_p <= Pix_119;
    10'd8:  neuron_3_mul_4_p <= Pix_120;
    10'd9:  neuron_3_mul_4_p <= Pix_121;
    10'd10:  neuron_3_mul_4_p <= Pix_122;
    10'd11:  neuron_3_mul_4_p <= Pix_123;
    10'd12:  neuron_3_mul_4_p <= Pix_124;
    10'd13:  neuron_3_mul_4_p <= Pix_125;
    10'd14:  neuron_3_mul_4_p <= Pix_126;
    10'd15:  neuron_3_mul_4_p <= Pix_127;
    10'd16:  neuron_3_mul_4_p <= Pix_128;
    10'd17:  neuron_3_mul_4_p <= Pix_129;
    10'd18:  neuron_3_mul_4_p <= Pix_130;
    10'd19:  neuron_3_mul_4_p <= Pix_131;
    10'd20:  neuron_3_mul_4_p <= Pix_132;
    10'd21:  neuron_3_mul_4_p <= Pix_133;
    10'd22:  neuron_3_mul_4_p <= Pix_134;
    10'd23:  neuron_3_mul_4_p <= Pix_135;
    10'd24:  neuron_3_mul_4_p <= Pix_136;
    10'd25:  neuron_3_mul_4_p <= Pix_137;
    10'd26:  neuron_3_mul_4_p <= Pix_138;
    10'd27:  neuron_3_mul_4_p <= Pix_139;
    default: neuron_3_mul_4_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_5_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_5_p <= Pix_140;
    10'd1:  neuron_3_mul_5_p <= Pix_141;
    10'd2:  neuron_3_mul_5_p <= Pix_142;
    10'd3:  neuron_3_mul_5_p <= Pix_143;
    10'd4:  neuron_3_mul_5_p <= Pix_144;
    10'd5:  neuron_3_mul_5_p <= Pix_145;
    10'd6:  neuron_3_mul_5_p <= Pix_146;
    10'd7:  neuron_3_mul_5_p <= Pix_147;
    10'd8:  neuron_3_mul_5_p <= Pix_148;
    10'd9:  neuron_3_mul_5_p <= Pix_149;
    10'd10:  neuron_3_mul_5_p <= Pix_150;
    10'd11:  neuron_3_mul_5_p <= Pix_151;
    10'd12:  neuron_3_mul_5_p <= Pix_152;
    10'd13:  neuron_3_mul_5_p <= Pix_153;
    10'd14:  neuron_3_mul_5_p <= Pix_154;
    10'd15:  neuron_3_mul_5_p <= Pix_155;
    10'd16:  neuron_3_mul_5_p <= Pix_156;
    10'd17:  neuron_3_mul_5_p <= Pix_157;
    10'd18:  neuron_3_mul_5_p <= Pix_158;
    10'd19:  neuron_3_mul_5_p <= Pix_159;
    10'd20:  neuron_3_mul_5_p <= Pix_160;
    10'd21:  neuron_3_mul_5_p <= Pix_161;
    10'd22:  neuron_3_mul_5_p <= Pix_162;
    10'd23:  neuron_3_mul_5_p <= Pix_163;
    10'd24:  neuron_3_mul_5_p <= Pix_164;
    10'd25:  neuron_3_mul_5_p <= Pix_165;
    10'd26:  neuron_3_mul_5_p <= Pix_166;
    10'd27:  neuron_3_mul_5_p <= Pix_167;
    default: neuron_3_mul_5_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_6_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_6_p <= Pix_168;
    10'd1:  neuron_3_mul_6_p <= Pix_169;
    10'd2:  neuron_3_mul_6_p <= Pix_170;
    10'd3:  neuron_3_mul_6_p <= Pix_171;
    10'd4:  neuron_3_mul_6_p <= Pix_172;
    10'd5:  neuron_3_mul_6_p <= Pix_173;
    10'd6:  neuron_3_mul_6_p <= Pix_174;
    10'd7:  neuron_3_mul_6_p <= Pix_175;
    10'd8:  neuron_3_mul_6_p <= Pix_176;
    10'd9:  neuron_3_mul_6_p <= Pix_177;
    10'd10:  neuron_3_mul_6_p <= Pix_178;
    10'd11:  neuron_3_mul_6_p <= Pix_179;
    10'd12:  neuron_3_mul_6_p <= Pix_180;
    10'd13:  neuron_3_mul_6_p <= Pix_181;
    10'd14:  neuron_3_mul_6_p <= Pix_182;
    10'd15:  neuron_3_mul_6_p <= Pix_183;
    10'd16:  neuron_3_mul_6_p <= Pix_184;
    10'd17:  neuron_3_mul_6_p <= Pix_185;
    10'd18:  neuron_3_mul_6_p <= Pix_186;
    10'd19:  neuron_3_mul_6_p <= Pix_187;
    10'd20:  neuron_3_mul_6_p <= Pix_188;
    10'd21:  neuron_3_mul_6_p <= Pix_189;
    10'd22:  neuron_3_mul_6_p <= Pix_190;
    10'd23:  neuron_3_mul_6_p <= Pix_191;
    10'd24:  neuron_3_mul_6_p <= Pix_192;
    10'd25:  neuron_3_mul_6_p <= Pix_193;
    10'd26:  neuron_3_mul_6_p <= Pix_194;
    10'd27:  neuron_3_mul_6_p <= Pix_195;
    default: neuron_3_mul_6_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_7_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_7_p <= Pix_196;
    10'd1:  neuron_3_mul_7_p <= Pix_197;
    10'd2:  neuron_3_mul_7_p <= Pix_198;
    10'd3:  neuron_3_mul_7_p <= Pix_199;
    10'd4:  neuron_3_mul_7_p <= Pix_200;
    10'd5:  neuron_3_mul_7_p <= Pix_201;
    10'd6:  neuron_3_mul_7_p <= Pix_202;
    10'd7:  neuron_3_mul_7_p <= Pix_203;
    10'd8:  neuron_3_mul_7_p <= Pix_204;
    10'd9:  neuron_3_mul_7_p <= Pix_205;
    10'd10:  neuron_3_mul_7_p <= Pix_206;
    10'd11:  neuron_3_mul_7_p <= Pix_207;
    10'd12:  neuron_3_mul_7_p <= Pix_208;
    10'd13:  neuron_3_mul_7_p <= Pix_209;
    10'd14:  neuron_3_mul_7_p <= Pix_210;
    10'd15:  neuron_3_mul_7_p <= Pix_211;
    10'd16:  neuron_3_mul_7_p <= Pix_212;
    10'd17:  neuron_3_mul_7_p <= Pix_213;
    10'd18:  neuron_3_mul_7_p <= Pix_214;
    10'd19:  neuron_3_mul_7_p <= Pix_215;
    10'd20:  neuron_3_mul_7_p <= Pix_216;
    10'd21:  neuron_3_mul_7_p <= Pix_217;
    10'd22:  neuron_3_mul_7_p <= Pix_218;
    10'd23:  neuron_3_mul_7_p <= Pix_219;
    10'd24:  neuron_3_mul_7_p <= Pix_220;
    10'd25:  neuron_3_mul_7_p <= Pix_221;
    10'd26:  neuron_3_mul_7_p <= Pix_222;
    10'd27:  neuron_3_mul_7_p <= Pix_223;
    default: neuron_3_mul_7_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_8_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_8_p <= Pix_224;
    10'd1:  neuron_3_mul_8_p <= Pix_225;
    10'd2:  neuron_3_mul_8_p <= Pix_226;
    10'd3:  neuron_3_mul_8_p <= Pix_227;
    10'd4:  neuron_3_mul_8_p <= Pix_228;
    10'd5:  neuron_3_mul_8_p <= Pix_229;
    10'd6:  neuron_3_mul_8_p <= Pix_230;
    10'd7:  neuron_3_mul_8_p <= Pix_231;
    10'd8:  neuron_3_mul_8_p <= Pix_232;
    10'd9:  neuron_3_mul_8_p <= Pix_233;
    10'd10:  neuron_3_mul_8_p <= Pix_234;
    10'd11:  neuron_3_mul_8_p <= Pix_235;
    10'd12:  neuron_3_mul_8_p <= Pix_236;
    10'd13:  neuron_3_mul_8_p <= Pix_237;
    10'd14:  neuron_3_mul_8_p <= Pix_238;
    10'd15:  neuron_3_mul_8_p <= Pix_239;
    10'd16:  neuron_3_mul_8_p <= Pix_240;
    10'd17:  neuron_3_mul_8_p <= Pix_241;
    10'd18:  neuron_3_mul_8_p <= Pix_242;
    10'd19:  neuron_3_mul_8_p <= Pix_243;
    10'd20:  neuron_3_mul_8_p <= Pix_244;
    10'd21:  neuron_3_mul_8_p <= Pix_245;
    10'd22:  neuron_3_mul_8_p <= Pix_246;
    10'd23:  neuron_3_mul_8_p <= Pix_247;
    10'd24:  neuron_3_mul_8_p <= Pix_248;
    10'd25:  neuron_3_mul_8_p <= Pix_249;
    10'd26:  neuron_3_mul_8_p <= Pix_250;
    10'd27:  neuron_3_mul_8_p <= Pix_251;
    default: neuron_3_mul_8_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_9_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_9_p <= Pix_252;
    10'd1:  neuron_3_mul_9_p <= Pix_253;
    10'd2:  neuron_3_mul_9_p <= Pix_254;
    10'd3:  neuron_3_mul_9_p <= Pix_255;
    10'd4:  neuron_3_mul_9_p <= Pix_256;
    10'd5:  neuron_3_mul_9_p <= Pix_257;
    10'd6:  neuron_3_mul_9_p <= Pix_258;
    10'd7:  neuron_3_mul_9_p <= Pix_259;
    10'd8:  neuron_3_mul_9_p <= Pix_260;
    10'd9:  neuron_3_mul_9_p <= Pix_261;
    10'd10:  neuron_3_mul_9_p <= Pix_262;
    10'd11:  neuron_3_mul_9_p <= Pix_263;
    10'd12:  neuron_3_mul_9_p <= Pix_264;
    10'd13:  neuron_3_mul_9_p <= Pix_265;
    10'd14:  neuron_3_mul_9_p <= Pix_266;
    10'd15:  neuron_3_mul_9_p <= Pix_267;
    10'd16:  neuron_3_mul_9_p <= Pix_268;
    10'd17:  neuron_3_mul_9_p <= Pix_269;
    10'd18:  neuron_3_mul_9_p <= Pix_270;
    10'd19:  neuron_3_mul_9_p <= Pix_271;
    10'd20:  neuron_3_mul_9_p <= Pix_272;
    10'd21:  neuron_3_mul_9_p <= Pix_273;
    10'd22:  neuron_3_mul_9_p <= Pix_274;
    10'd23:  neuron_3_mul_9_p <= Pix_275;
    10'd24:  neuron_3_mul_9_p <= Pix_276;
    10'd25:  neuron_3_mul_9_p <= Pix_277;
    10'd26:  neuron_3_mul_9_p <= Pix_278;
    10'd27:  neuron_3_mul_9_p <= Pix_279;
    default: neuron_3_mul_9_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_10_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_10_p <= Pix_280;
    10'd1:  neuron_3_mul_10_p <= Pix_281;
    10'd2:  neuron_3_mul_10_p <= Pix_282;
    10'd3:  neuron_3_mul_10_p <= Pix_283;
    10'd4:  neuron_3_mul_10_p <= Pix_284;
    10'd5:  neuron_3_mul_10_p <= Pix_285;
    10'd6:  neuron_3_mul_10_p <= Pix_286;
    10'd7:  neuron_3_mul_10_p <= Pix_287;
    10'd8:  neuron_3_mul_10_p <= Pix_288;
    10'd9:  neuron_3_mul_10_p <= Pix_289;
    10'd10:  neuron_3_mul_10_p <= Pix_290;
    10'd11:  neuron_3_mul_10_p <= Pix_291;
    10'd12:  neuron_3_mul_10_p <= Pix_292;
    10'd13:  neuron_3_mul_10_p <= Pix_293;
    10'd14:  neuron_3_mul_10_p <= Pix_294;
    10'd15:  neuron_3_mul_10_p <= Pix_295;
    10'd16:  neuron_3_mul_10_p <= Pix_296;
    10'd17:  neuron_3_mul_10_p <= Pix_297;
    10'd18:  neuron_3_mul_10_p <= Pix_298;
    10'd19:  neuron_3_mul_10_p <= Pix_299;
    10'd20:  neuron_3_mul_10_p <= Pix_300;
    10'd21:  neuron_3_mul_10_p <= Pix_301;
    10'd22:  neuron_3_mul_10_p <= Pix_302;
    10'd23:  neuron_3_mul_10_p <= Pix_303;
    10'd24:  neuron_3_mul_10_p <= Pix_304;
    10'd25:  neuron_3_mul_10_p <= Pix_305;
    10'd26:  neuron_3_mul_10_p <= Pix_306;
    10'd27:  neuron_3_mul_10_p <= Pix_307;
    default: neuron_3_mul_10_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_11_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_11_p <= Pix_308;
    10'd1:  neuron_3_mul_11_p <= Pix_309;
    10'd2:  neuron_3_mul_11_p <= Pix_310;
    10'd3:  neuron_3_mul_11_p <= Pix_311;
    10'd4:  neuron_3_mul_11_p <= Pix_312;
    10'd5:  neuron_3_mul_11_p <= Pix_313;
    10'd6:  neuron_3_mul_11_p <= Pix_314;
    10'd7:  neuron_3_mul_11_p <= Pix_315;
    10'd8:  neuron_3_mul_11_p <= Pix_316;
    10'd9:  neuron_3_mul_11_p <= Pix_317;
    10'd10:  neuron_3_mul_11_p <= Pix_318;
    10'd11:  neuron_3_mul_11_p <= Pix_319;
    10'd12:  neuron_3_mul_11_p <= Pix_320;
    10'd13:  neuron_3_mul_11_p <= Pix_321;
    10'd14:  neuron_3_mul_11_p <= Pix_322;
    10'd15:  neuron_3_mul_11_p <= Pix_323;
    10'd16:  neuron_3_mul_11_p <= Pix_324;
    10'd17:  neuron_3_mul_11_p <= Pix_325;
    10'd18:  neuron_3_mul_11_p <= Pix_326;
    10'd19:  neuron_3_mul_11_p <= Pix_327;
    10'd20:  neuron_3_mul_11_p <= Pix_328;
    10'd21:  neuron_3_mul_11_p <= Pix_329;
    10'd22:  neuron_3_mul_11_p <= Pix_330;
    10'd23:  neuron_3_mul_11_p <= Pix_331;
    10'd24:  neuron_3_mul_11_p <= Pix_332;
    10'd25:  neuron_3_mul_11_p <= Pix_333;
    10'd26:  neuron_3_mul_11_p <= Pix_334;
    10'd27:  neuron_3_mul_11_p <= Pix_335;
    default: neuron_3_mul_11_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_12_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_12_p <= Pix_336;
    10'd1:  neuron_3_mul_12_p <= Pix_337;
    10'd2:  neuron_3_mul_12_p <= Pix_338;
    10'd3:  neuron_3_mul_12_p <= Pix_339;
    10'd4:  neuron_3_mul_12_p <= Pix_340;
    10'd5:  neuron_3_mul_12_p <= Pix_341;
    10'd6:  neuron_3_mul_12_p <= Pix_342;
    10'd7:  neuron_3_mul_12_p <= Pix_343;
    10'd8:  neuron_3_mul_12_p <= Pix_344;
    10'd9:  neuron_3_mul_12_p <= Pix_345;
    10'd10:  neuron_3_mul_12_p <= Pix_346;
    10'd11:  neuron_3_mul_12_p <= Pix_347;
    10'd12:  neuron_3_mul_12_p <= Pix_348;
    10'd13:  neuron_3_mul_12_p <= Pix_349;
    10'd14:  neuron_3_mul_12_p <= Pix_350;
    10'd15:  neuron_3_mul_12_p <= Pix_351;
    10'd16:  neuron_3_mul_12_p <= Pix_352;
    10'd17:  neuron_3_mul_12_p <= Pix_353;
    10'd18:  neuron_3_mul_12_p <= Pix_354;
    10'd19:  neuron_3_mul_12_p <= Pix_355;
    10'd20:  neuron_3_mul_12_p <= Pix_356;
    10'd21:  neuron_3_mul_12_p <= Pix_357;
    10'd22:  neuron_3_mul_12_p <= Pix_358;
    10'd23:  neuron_3_mul_12_p <= Pix_359;
    10'd24:  neuron_3_mul_12_p <= Pix_360;
    10'd25:  neuron_3_mul_12_p <= Pix_361;
    10'd26:  neuron_3_mul_12_p <= Pix_362;
    10'd27:  neuron_3_mul_12_p <= Pix_363;
    default: neuron_3_mul_12_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_13_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_13_p <= Pix_364;
    10'd1:  neuron_3_mul_13_p <= Pix_365;
    10'd2:  neuron_3_mul_13_p <= Pix_366;
    10'd3:  neuron_3_mul_13_p <= Pix_367;
    10'd4:  neuron_3_mul_13_p <= Pix_368;
    10'd5:  neuron_3_mul_13_p <= Pix_369;
    10'd6:  neuron_3_mul_13_p <= Pix_370;
    10'd7:  neuron_3_mul_13_p <= Pix_371;
    10'd8:  neuron_3_mul_13_p <= Pix_372;
    10'd9:  neuron_3_mul_13_p <= Pix_373;
    10'd10:  neuron_3_mul_13_p <= Pix_374;
    10'd11:  neuron_3_mul_13_p <= Pix_375;
    10'd12:  neuron_3_mul_13_p <= Pix_376;
    10'd13:  neuron_3_mul_13_p <= Pix_377;
    10'd14:  neuron_3_mul_13_p <= Pix_378;
    10'd15:  neuron_3_mul_13_p <= Pix_379;
    10'd16:  neuron_3_mul_13_p <= Pix_380;
    10'd17:  neuron_3_mul_13_p <= Pix_381;
    10'd18:  neuron_3_mul_13_p <= Pix_382;
    10'd19:  neuron_3_mul_13_p <= Pix_383;
    10'd20:  neuron_3_mul_13_p <= Pix_384;
    10'd21:  neuron_3_mul_13_p <= Pix_385;
    10'd22:  neuron_3_mul_13_p <= Pix_386;
    10'd23:  neuron_3_mul_13_p <= Pix_387;
    10'd24:  neuron_3_mul_13_p <= Pix_388;
    10'd25:  neuron_3_mul_13_p <= Pix_389;
    10'd26:  neuron_3_mul_13_p <= Pix_390;
    10'd27:  neuron_3_mul_13_p <= Pix_391;
    default: neuron_3_mul_13_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_14_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_14_p <= Pix_392;
    10'd1:  neuron_3_mul_14_p <= Pix_393;
    10'd2:  neuron_3_mul_14_p <= Pix_394;
    10'd3:  neuron_3_mul_14_p <= Pix_395;
    10'd4:  neuron_3_mul_14_p <= Pix_396;
    10'd5:  neuron_3_mul_14_p <= Pix_397;
    10'd6:  neuron_3_mul_14_p <= Pix_398;
    10'd7:  neuron_3_mul_14_p <= Pix_399;
    10'd8:  neuron_3_mul_14_p <= Pix_400;
    10'd9:  neuron_3_mul_14_p <= Pix_401;
    10'd10:  neuron_3_mul_14_p <= Pix_402;
    10'd11:  neuron_3_mul_14_p <= Pix_403;
    10'd12:  neuron_3_mul_14_p <= Pix_404;
    10'd13:  neuron_3_mul_14_p <= Pix_405;
    10'd14:  neuron_3_mul_14_p <= Pix_406;
    10'd15:  neuron_3_mul_14_p <= Pix_407;
    10'd16:  neuron_3_mul_14_p <= Pix_408;
    10'd17:  neuron_3_mul_14_p <= Pix_409;
    10'd18:  neuron_3_mul_14_p <= Pix_410;
    10'd19:  neuron_3_mul_14_p <= Pix_411;
    10'd20:  neuron_3_mul_14_p <= Pix_412;
    10'd21:  neuron_3_mul_14_p <= Pix_413;
    10'd22:  neuron_3_mul_14_p <= Pix_414;
    10'd23:  neuron_3_mul_14_p <= Pix_415;
    10'd24:  neuron_3_mul_14_p <= Pix_416;
    10'd25:  neuron_3_mul_14_p <= Pix_417;
    10'd26:  neuron_3_mul_14_p <= Pix_418;
    10'd27:  neuron_3_mul_14_p <= Pix_419;
    default: neuron_3_mul_14_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_15_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_15_p <= Pix_420;
    10'd1:  neuron_3_mul_15_p <= Pix_421;
    10'd2:  neuron_3_mul_15_p <= Pix_422;
    10'd3:  neuron_3_mul_15_p <= Pix_423;
    10'd4:  neuron_3_mul_15_p <= Pix_424;
    10'd5:  neuron_3_mul_15_p <= Pix_425;
    10'd6:  neuron_3_mul_15_p <= Pix_426;
    10'd7:  neuron_3_mul_15_p <= Pix_427;
    10'd8:  neuron_3_mul_15_p <= Pix_428;
    10'd9:  neuron_3_mul_15_p <= Pix_429;
    10'd10:  neuron_3_mul_15_p <= Pix_430;
    10'd11:  neuron_3_mul_15_p <= Pix_431;
    10'd12:  neuron_3_mul_15_p <= Pix_432;
    10'd13:  neuron_3_mul_15_p <= Pix_433;
    10'd14:  neuron_3_mul_15_p <= Pix_434;
    10'd15:  neuron_3_mul_15_p <= Pix_435;
    10'd16:  neuron_3_mul_15_p <= Pix_436;
    10'd17:  neuron_3_mul_15_p <= Pix_437;
    10'd18:  neuron_3_mul_15_p <= Pix_438;
    10'd19:  neuron_3_mul_15_p <= Pix_439;
    10'd20:  neuron_3_mul_15_p <= Pix_440;
    10'd21:  neuron_3_mul_15_p <= Pix_441;
    10'd22:  neuron_3_mul_15_p <= Pix_442;
    10'd23:  neuron_3_mul_15_p <= Pix_443;
    10'd24:  neuron_3_mul_15_p <= Pix_444;
    10'd25:  neuron_3_mul_15_p <= Pix_445;
    10'd26:  neuron_3_mul_15_p <= Pix_446;
    10'd27:  neuron_3_mul_15_p <= Pix_447;
    default: neuron_3_mul_15_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_16_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_16_p <= Pix_448;
    10'd1:  neuron_3_mul_16_p <= Pix_449;
    10'd2:  neuron_3_mul_16_p <= Pix_450;
    10'd3:  neuron_3_mul_16_p <= Pix_451;
    10'd4:  neuron_3_mul_16_p <= Pix_452;
    10'd5:  neuron_3_mul_16_p <= Pix_453;
    10'd6:  neuron_3_mul_16_p <= Pix_454;
    10'd7:  neuron_3_mul_16_p <= Pix_455;
    10'd8:  neuron_3_mul_16_p <= Pix_456;
    10'd9:  neuron_3_mul_16_p <= Pix_457;
    10'd10:  neuron_3_mul_16_p <= Pix_458;
    10'd11:  neuron_3_mul_16_p <= Pix_459;
    10'd12:  neuron_3_mul_16_p <= Pix_460;
    10'd13:  neuron_3_mul_16_p <= Pix_461;
    10'd14:  neuron_3_mul_16_p <= Pix_462;
    10'd15:  neuron_3_mul_16_p <= Pix_463;
    10'd16:  neuron_3_mul_16_p <= Pix_464;
    10'd17:  neuron_3_mul_16_p <= Pix_465;
    10'd18:  neuron_3_mul_16_p <= Pix_466;
    10'd19:  neuron_3_mul_16_p <= Pix_467;
    10'd20:  neuron_3_mul_16_p <= Pix_468;
    10'd21:  neuron_3_mul_16_p <= Pix_469;
    10'd22:  neuron_3_mul_16_p <= Pix_470;
    10'd23:  neuron_3_mul_16_p <= Pix_471;
    10'd24:  neuron_3_mul_16_p <= Pix_472;
    10'd25:  neuron_3_mul_16_p <= Pix_473;
    10'd26:  neuron_3_mul_16_p <= Pix_474;
    10'd27:  neuron_3_mul_16_p <= Pix_475;
    default: neuron_3_mul_16_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_17_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_17_p <= Pix_476;
    10'd1:  neuron_3_mul_17_p <= Pix_477;
    10'd2:  neuron_3_mul_17_p <= Pix_478;
    10'd3:  neuron_3_mul_17_p <= Pix_479;
    10'd4:  neuron_3_mul_17_p <= Pix_480;
    10'd5:  neuron_3_mul_17_p <= Pix_481;
    10'd6:  neuron_3_mul_17_p <= Pix_482;
    10'd7:  neuron_3_mul_17_p <= Pix_483;
    10'd8:  neuron_3_mul_17_p <= Pix_484;
    10'd9:  neuron_3_mul_17_p <= Pix_485;
    10'd10:  neuron_3_mul_17_p <= Pix_486;
    10'd11:  neuron_3_mul_17_p <= Pix_487;
    10'd12:  neuron_3_mul_17_p <= Pix_488;
    10'd13:  neuron_3_mul_17_p <= Pix_489;
    10'd14:  neuron_3_mul_17_p <= Pix_490;
    10'd15:  neuron_3_mul_17_p <= Pix_491;
    10'd16:  neuron_3_mul_17_p <= Pix_492;
    10'd17:  neuron_3_mul_17_p <= Pix_493;
    10'd18:  neuron_3_mul_17_p <= Pix_494;
    10'd19:  neuron_3_mul_17_p <= Pix_495;
    10'd20:  neuron_3_mul_17_p <= Pix_496;
    10'd21:  neuron_3_mul_17_p <= Pix_497;
    10'd22:  neuron_3_mul_17_p <= Pix_498;
    10'd23:  neuron_3_mul_17_p <= Pix_499;
    10'd24:  neuron_3_mul_17_p <= Pix_500;
    10'd25:  neuron_3_mul_17_p <= Pix_501;
    10'd26:  neuron_3_mul_17_p <= Pix_502;
    10'd27:  neuron_3_mul_17_p <= Pix_503;
    default: neuron_3_mul_17_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_18_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_18_p <= Pix_504;
    10'd1:  neuron_3_mul_18_p <= Pix_505;
    10'd2:  neuron_3_mul_18_p <= Pix_506;
    10'd3:  neuron_3_mul_18_p <= Pix_507;
    10'd4:  neuron_3_mul_18_p <= Pix_508;
    10'd5:  neuron_3_mul_18_p <= Pix_509;
    10'd6:  neuron_3_mul_18_p <= Pix_510;
    10'd7:  neuron_3_mul_18_p <= Pix_511;
    10'd8:  neuron_3_mul_18_p <= Pix_512;
    10'd9:  neuron_3_mul_18_p <= Pix_513;
    10'd10:  neuron_3_mul_18_p <= Pix_514;
    10'd11:  neuron_3_mul_18_p <= Pix_515;
    10'd12:  neuron_3_mul_18_p <= Pix_516;
    10'd13:  neuron_3_mul_18_p <= Pix_517;
    10'd14:  neuron_3_mul_18_p <= Pix_518;
    10'd15:  neuron_3_mul_18_p <= Pix_519;
    10'd16:  neuron_3_mul_18_p <= Pix_520;
    10'd17:  neuron_3_mul_18_p <= Pix_521;
    10'd18:  neuron_3_mul_18_p <= Pix_522;
    10'd19:  neuron_3_mul_18_p <= Pix_523;
    10'd20:  neuron_3_mul_18_p <= Pix_524;
    10'd21:  neuron_3_mul_18_p <= Pix_525;
    10'd22:  neuron_3_mul_18_p <= Pix_526;
    10'd23:  neuron_3_mul_18_p <= Pix_527;
    10'd24:  neuron_3_mul_18_p <= Pix_528;
    10'd25:  neuron_3_mul_18_p <= Pix_529;
    10'd26:  neuron_3_mul_18_p <= Pix_530;
    10'd27:  neuron_3_mul_18_p <= Pix_531;
    default: neuron_3_mul_18_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_19_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_19_p <= Pix_532;
    10'd1:  neuron_3_mul_19_p <= Pix_533;
    10'd2:  neuron_3_mul_19_p <= Pix_534;
    10'd3:  neuron_3_mul_19_p <= Pix_535;
    10'd4:  neuron_3_mul_19_p <= Pix_536;
    10'd5:  neuron_3_mul_19_p <= Pix_537;
    10'd6:  neuron_3_mul_19_p <= Pix_538;
    10'd7:  neuron_3_mul_19_p <= Pix_539;
    10'd8:  neuron_3_mul_19_p <= Pix_540;
    10'd9:  neuron_3_mul_19_p <= Pix_541;
    10'd10:  neuron_3_mul_19_p <= Pix_542;
    10'd11:  neuron_3_mul_19_p <= Pix_543;
    10'd12:  neuron_3_mul_19_p <= Pix_544;
    10'd13:  neuron_3_mul_19_p <= Pix_545;
    10'd14:  neuron_3_mul_19_p <= Pix_546;
    10'd15:  neuron_3_mul_19_p <= Pix_547;
    10'd16:  neuron_3_mul_19_p <= Pix_548;
    10'd17:  neuron_3_mul_19_p <= Pix_549;
    10'd18:  neuron_3_mul_19_p <= Pix_550;
    10'd19:  neuron_3_mul_19_p <= Pix_551;
    10'd20:  neuron_3_mul_19_p <= Pix_552;
    10'd21:  neuron_3_mul_19_p <= Pix_553;
    10'd22:  neuron_3_mul_19_p <= Pix_554;
    10'd23:  neuron_3_mul_19_p <= Pix_555;
    10'd24:  neuron_3_mul_19_p <= Pix_556;
    10'd25:  neuron_3_mul_19_p <= Pix_557;
    10'd26:  neuron_3_mul_19_p <= Pix_558;
    10'd27:  neuron_3_mul_19_p <= Pix_559;
    default: neuron_3_mul_19_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_20_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_20_p <= Pix_560;
    10'd1:  neuron_3_mul_20_p <= Pix_561;
    10'd2:  neuron_3_mul_20_p <= Pix_562;
    10'd3:  neuron_3_mul_20_p <= Pix_563;
    10'd4:  neuron_3_mul_20_p <= Pix_564;
    10'd5:  neuron_3_mul_20_p <= Pix_565;
    10'd6:  neuron_3_mul_20_p <= Pix_566;
    10'd7:  neuron_3_mul_20_p <= Pix_567;
    10'd8:  neuron_3_mul_20_p <= Pix_568;
    10'd9:  neuron_3_mul_20_p <= Pix_569;
    10'd10:  neuron_3_mul_20_p <= Pix_570;
    10'd11:  neuron_3_mul_20_p <= Pix_571;
    10'd12:  neuron_3_mul_20_p <= Pix_572;
    10'd13:  neuron_3_mul_20_p <= Pix_573;
    10'd14:  neuron_3_mul_20_p <= Pix_574;
    10'd15:  neuron_3_mul_20_p <= Pix_575;
    10'd16:  neuron_3_mul_20_p <= Pix_576;
    10'd17:  neuron_3_mul_20_p <= Pix_577;
    10'd18:  neuron_3_mul_20_p <= Pix_578;
    10'd19:  neuron_3_mul_20_p <= Pix_579;
    10'd20:  neuron_3_mul_20_p <= Pix_580;
    10'd21:  neuron_3_mul_20_p <= Pix_581;
    10'd22:  neuron_3_mul_20_p <= Pix_582;
    10'd23:  neuron_3_mul_20_p <= Pix_583;
    10'd24:  neuron_3_mul_20_p <= Pix_584;
    10'd25:  neuron_3_mul_20_p <= Pix_585;
    10'd26:  neuron_3_mul_20_p <= Pix_586;
    10'd27:  neuron_3_mul_20_p <= Pix_587;
    default: neuron_3_mul_20_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_21_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_21_p <= Pix_588;
    10'd1:  neuron_3_mul_21_p <= Pix_589;
    10'd2:  neuron_3_mul_21_p <= Pix_590;
    10'd3:  neuron_3_mul_21_p <= Pix_591;
    10'd4:  neuron_3_mul_21_p <= Pix_592;
    10'd5:  neuron_3_mul_21_p <= Pix_593;
    10'd6:  neuron_3_mul_21_p <= Pix_594;
    10'd7:  neuron_3_mul_21_p <= Pix_595;
    10'd8:  neuron_3_mul_21_p <= Pix_596;
    10'd9:  neuron_3_mul_21_p <= Pix_597;
    10'd10:  neuron_3_mul_21_p <= Pix_598;
    10'd11:  neuron_3_mul_21_p <= Pix_599;
    10'd12:  neuron_3_mul_21_p <= Pix_600;
    10'd13:  neuron_3_mul_21_p <= Pix_601;
    10'd14:  neuron_3_mul_21_p <= Pix_602;
    10'd15:  neuron_3_mul_21_p <= Pix_603;
    10'd16:  neuron_3_mul_21_p <= Pix_604;
    10'd17:  neuron_3_mul_21_p <= Pix_605;
    10'd18:  neuron_3_mul_21_p <= Pix_606;
    10'd19:  neuron_3_mul_21_p <= Pix_607;
    10'd20:  neuron_3_mul_21_p <= Pix_608;
    10'd21:  neuron_3_mul_21_p <= Pix_609;
    10'd22:  neuron_3_mul_21_p <= Pix_610;
    10'd23:  neuron_3_mul_21_p <= Pix_611;
    10'd24:  neuron_3_mul_21_p <= Pix_612;
    10'd25:  neuron_3_mul_21_p <= Pix_613;
    10'd26:  neuron_3_mul_21_p <= Pix_614;
    10'd27:  neuron_3_mul_21_p <= Pix_615;
    default: neuron_3_mul_21_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_22_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_22_p <= Pix_616;
    10'd1:  neuron_3_mul_22_p <= Pix_617;
    10'd2:  neuron_3_mul_22_p <= Pix_618;
    10'd3:  neuron_3_mul_22_p <= Pix_619;
    10'd4:  neuron_3_mul_22_p <= Pix_620;
    10'd5:  neuron_3_mul_22_p <= Pix_621;
    10'd6:  neuron_3_mul_22_p <= Pix_622;
    10'd7:  neuron_3_mul_22_p <= Pix_623;
    10'd8:  neuron_3_mul_22_p <= Pix_624;
    10'd9:  neuron_3_mul_22_p <= Pix_625;
    10'd10:  neuron_3_mul_22_p <= Pix_626;
    10'd11:  neuron_3_mul_22_p <= Pix_627;
    10'd12:  neuron_3_mul_22_p <= Pix_628;
    10'd13:  neuron_3_mul_22_p <= Pix_629;
    10'd14:  neuron_3_mul_22_p <= Pix_630;
    10'd15:  neuron_3_mul_22_p <= Pix_631;
    10'd16:  neuron_3_mul_22_p <= Pix_632;
    10'd17:  neuron_3_mul_22_p <= Pix_633;
    10'd18:  neuron_3_mul_22_p <= Pix_634;
    10'd19:  neuron_3_mul_22_p <= Pix_635;
    10'd20:  neuron_3_mul_22_p <= Pix_636;
    10'd21:  neuron_3_mul_22_p <= Pix_637;
    10'd22:  neuron_3_mul_22_p <= Pix_638;
    10'd23:  neuron_3_mul_22_p <= Pix_639;
    10'd24:  neuron_3_mul_22_p <= Pix_640;
    10'd25:  neuron_3_mul_22_p <= Pix_641;
    10'd26:  neuron_3_mul_22_p <= Pix_642;
    10'd27:  neuron_3_mul_22_p <= Pix_643;
    default: neuron_3_mul_22_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_23_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_23_p <= Pix_644;
    10'd1:  neuron_3_mul_23_p <= Pix_645;
    10'd2:  neuron_3_mul_23_p <= Pix_646;
    10'd3:  neuron_3_mul_23_p <= Pix_647;
    10'd4:  neuron_3_mul_23_p <= Pix_648;
    10'd5:  neuron_3_mul_23_p <= Pix_649;
    10'd6:  neuron_3_mul_23_p <= Pix_650;
    10'd7:  neuron_3_mul_23_p <= Pix_651;
    10'd8:  neuron_3_mul_23_p <= Pix_652;
    10'd9:  neuron_3_mul_23_p <= Pix_653;
    10'd10:  neuron_3_mul_23_p <= Pix_654;
    10'd11:  neuron_3_mul_23_p <= Pix_655;
    10'd12:  neuron_3_mul_23_p <= Pix_656;
    10'd13:  neuron_3_mul_23_p <= Pix_657;
    10'd14:  neuron_3_mul_23_p <= Pix_658;
    10'd15:  neuron_3_mul_23_p <= Pix_659;
    10'd16:  neuron_3_mul_23_p <= Pix_660;
    10'd17:  neuron_3_mul_23_p <= Pix_661;
    10'd18:  neuron_3_mul_23_p <= Pix_662;
    10'd19:  neuron_3_mul_23_p <= Pix_663;
    10'd20:  neuron_3_mul_23_p <= Pix_664;
    10'd21:  neuron_3_mul_23_p <= Pix_665;
    10'd22:  neuron_3_mul_23_p <= Pix_666;
    10'd23:  neuron_3_mul_23_p <= Pix_667;
    10'd24:  neuron_3_mul_23_p <= Pix_668;
    10'd25:  neuron_3_mul_23_p <= Pix_669;
    10'd26:  neuron_3_mul_23_p <= Pix_670;
    10'd27:  neuron_3_mul_23_p <= Pix_671;
    default: neuron_3_mul_23_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_24_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_24_p <= Pix_672;
    10'd1:  neuron_3_mul_24_p <= Pix_673;
    10'd2:  neuron_3_mul_24_p <= Pix_674;
    10'd3:  neuron_3_mul_24_p <= Pix_675;
    10'd4:  neuron_3_mul_24_p <= Pix_676;
    10'd5:  neuron_3_mul_24_p <= Pix_677;
    10'd6:  neuron_3_mul_24_p <= Pix_678;
    10'd7:  neuron_3_mul_24_p <= Pix_679;
    10'd8:  neuron_3_mul_24_p <= Pix_680;
    10'd9:  neuron_3_mul_24_p <= Pix_681;
    10'd10:  neuron_3_mul_24_p <= Pix_682;
    10'd11:  neuron_3_mul_24_p <= Pix_683;
    10'd12:  neuron_3_mul_24_p <= Pix_684;
    10'd13:  neuron_3_mul_24_p <= Pix_685;
    10'd14:  neuron_3_mul_24_p <= Pix_686;
    10'd15:  neuron_3_mul_24_p <= Pix_687;
    10'd16:  neuron_3_mul_24_p <= Pix_688;
    10'd17:  neuron_3_mul_24_p <= Pix_689;
    10'd18:  neuron_3_mul_24_p <= Pix_690;
    10'd19:  neuron_3_mul_24_p <= Pix_691;
    10'd20:  neuron_3_mul_24_p <= Pix_692;
    10'd21:  neuron_3_mul_24_p <= Pix_693;
    10'd22:  neuron_3_mul_24_p <= Pix_694;
    10'd23:  neuron_3_mul_24_p <= Pix_695;
    10'd24:  neuron_3_mul_24_p <= Pix_696;
    10'd25:  neuron_3_mul_24_p <= Pix_697;
    10'd26:  neuron_3_mul_24_p <= Pix_698;
    10'd27:  neuron_3_mul_24_p <= Pix_699;
    default: neuron_3_mul_24_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_25_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_25_p <= Pix_700;
    10'd1:  neuron_3_mul_25_p <= Pix_701;
    10'd2:  neuron_3_mul_25_p <= Pix_702;
    10'd3:  neuron_3_mul_25_p <= Pix_703;
    10'd4:  neuron_3_mul_25_p <= Pix_704;
    10'd5:  neuron_3_mul_25_p <= Pix_705;
    10'd6:  neuron_3_mul_25_p <= Pix_706;
    10'd7:  neuron_3_mul_25_p <= Pix_707;
    10'd8:  neuron_3_mul_25_p <= Pix_708;
    10'd9:  neuron_3_mul_25_p <= Pix_709;
    10'd10:  neuron_3_mul_25_p <= Pix_710;
    10'd11:  neuron_3_mul_25_p <= Pix_711;
    10'd12:  neuron_3_mul_25_p <= Pix_712;
    10'd13:  neuron_3_mul_25_p <= Pix_713;
    10'd14:  neuron_3_mul_25_p <= Pix_714;
    10'd15:  neuron_3_mul_25_p <= Pix_715;
    10'd16:  neuron_3_mul_25_p <= Pix_716;
    10'd17:  neuron_3_mul_25_p <= Pix_717;
    10'd18:  neuron_3_mul_25_p <= Pix_718;
    10'd19:  neuron_3_mul_25_p <= Pix_719;
    10'd20:  neuron_3_mul_25_p <= Pix_720;
    10'd21:  neuron_3_mul_25_p <= Pix_721;
    10'd22:  neuron_3_mul_25_p <= Pix_722;
    10'd23:  neuron_3_mul_25_p <= Pix_723;
    10'd24:  neuron_3_mul_25_p <= Pix_724;
    10'd25:  neuron_3_mul_25_p <= Pix_725;
    10'd26:  neuron_3_mul_25_p <= Pix_726;
    10'd27:  neuron_3_mul_25_p <= Pix_727;
    default: neuron_3_mul_25_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_26_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_26_p <= Pix_728;
    10'd1:  neuron_3_mul_26_p <= Pix_729;
    10'd2:  neuron_3_mul_26_p <= Pix_730;
    10'd3:  neuron_3_mul_26_p <= Pix_731;
    10'd4:  neuron_3_mul_26_p <= Pix_732;
    10'd5:  neuron_3_mul_26_p <= Pix_733;
    10'd6:  neuron_3_mul_26_p <= Pix_734;
    10'd7:  neuron_3_mul_26_p <= Pix_735;
    10'd8:  neuron_3_mul_26_p <= Pix_736;
    10'd9:  neuron_3_mul_26_p <= Pix_737;
    10'd10:  neuron_3_mul_26_p <= Pix_738;
    10'd11:  neuron_3_mul_26_p <= Pix_739;
    10'd12:  neuron_3_mul_26_p <= Pix_740;
    10'd13:  neuron_3_mul_26_p <= Pix_741;
    10'd14:  neuron_3_mul_26_p <= Pix_742;
    10'd15:  neuron_3_mul_26_p <= Pix_743;
    10'd16:  neuron_3_mul_26_p <= Pix_744;
    10'd17:  neuron_3_mul_26_p <= Pix_745;
    10'd18:  neuron_3_mul_26_p <= Pix_746;
    10'd19:  neuron_3_mul_26_p <= Pix_747;
    10'd20:  neuron_3_mul_26_p <= Pix_748;
    10'd21:  neuron_3_mul_26_p <= Pix_749;
    10'd22:  neuron_3_mul_26_p <= Pix_750;
    10'd23:  neuron_3_mul_26_p <= Pix_751;
    10'd24:  neuron_3_mul_26_p <= Pix_752;
    10'd25:  neuron_3_mul_26_p <= Pix_753;
    10'd26:  neuron_3_mul_26_p <= Pix_754;
    10'd27:  neuron_3_mul_26_p <= Pix_755;
    default: neuron_3_mul_26_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_3_mul_27_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_3_mul_27_p <= Pix_756;
    10'd1:  neuron_3_mul_27_p <= Pix_757;
    10'd2:  neuron_3_mul_27_p <= Pix_758;
    10'd3:  neuron_3_mul_27_p <= Pix_759;
    10'd4:  neuron_3_mul_27_p <= Pix_760;
    10'd5:  neuron_3_mul_27_p <= Pix_761;
    10'd6:  neuron_3_mul_27_p <= Pix_762;
    10'd7:  neuron_3_mul_27_p <= Pix_763;
    10'd8:  neuron_3_mul_27_p <= Pix_764;
    10'd9:  neuron_3_mul_27_p <= Pix_765;
    10'd10:  neuron_3_mul_27_p <= Pix_766;
    10'd11:  neuron_3_mul_27_p <= Pix_767;
    10'd12:  neuron_3_mul_27_p <= Pix_768;
    10'd13:  neuron_3_mul_27_p <= Pix_769;
    10'd14:  neuron_3_mul_27_p <= Pix_770;
    10'd15:  neuron_3_mul_27_p <= Pix_771;
    10'd16:  neuron_3_mul_27_p <= Pix_772;
    10'd17:  neuron_3_mul_27_p <= Pix_773;
    10'd18:  neuron_3_mul_27_p <= Pix_774;
    10'd19:  neuron_3_mul_27_p <= Pix_775;
    10'd20:  neuron_3_mul_27_p <= Pix_776;
    10'd21:  neuron_3_mul_27_p <= Pix_777;
    10'd22:  neuron_3_mul_27_p <= Pix_778;
    10'd23:  neuron_3_mul_27_p <= Pix_779;
    10'd24:  neuron_3_mul_27_p <= Pix_780;
    10'd25:  neuron_3_mul_27_p <= Pix_781;
    10'd26:  neuron_3_mul_27_p <= Pix_782;
    10'd27:  neuron_3_mul_27_p <= Pix_783;
    default: neuron_3_mul_27_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_0_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_0_p <= Pix_0;
    10'd1:  neuron_4_mul_0_p <= Pix_1;
    10'd2:  neuron_4_mul_0_p <= Pix_2;
    10'd3:  neuron_4_mul_0_p <= Pix_3;
    10'd4:  neuron_4_mul_0_p <= Pix_4;
    10'd5:  neuron_4_mul_0_p <= Pix_5;
    10'd6:  neuron_4_mul_0_p <= Pix_6;
    10'd7:  neuron_4_mul_0_p <= Pix_7;
    10'd8:  neuron_4_mul_0_p <= Pix_8;
    10'd9:  neuron_4_mul_0_p <= Pix_9;
    10'd10:  neuron_4_mul_0_p <= Pix_10;
    10'd11:  neuron_4_mul_0_p <= Pix_11;
    10'd12:  neuron_4_mul_0_p <= Pix_12;
    10'd13:  neuron_4_mul_0_p <= Pix_13;
    10'd14:  neuron_4_mul_0_p <= Pix_14;
    10'd15:  neuron_4_mul_0_p <= Pix_15;
    10'd16:  neuron_4_mul_0_p <= Pix_16;
    10'd17:  neuron_4_mul_0_p <= Pix_17;
    10'd18:  neuron_4_mul_0_p <= Pix_18;
    10'd19:  neuron_4_mul_0_p <= Pix_19;
    10'd20:  neuron_4_mul_0_p <= Pix_20;
    10'd21:  neuron_4_mul_0_p <= Pix_21;
    10'd22:  neuron_4_mul_0_p <= Pix_22;
    10'd23:  neuron_4_mul_0_p <= Pix_23;
    10'd24:  neuron_4_mul_0_p <= Pix_24;
    10'd25:  neuron_4_mul_0_p <= Pix_25;
    10'd26:  neuron_4_mul_0_p <= Pix_26;
    10'd27:  neuron_4_mul_0_p <= Pix_27;
    default: neuron_4_mul_0_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_1_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_1_p <= Pix_28;
    10'd1:  neuron_4_mul_1_p <= Pix_29;
    10'd2:  neuron_4_mul_1_p <= Pix_30;
    10'd3:  neuron_4_mul_1_p <= Pix_31;
    10'd4:  neuron_4_mul_1_p <= Pix_32;
    10'd5:  neuron_4_mul_1_p <= Pix_33;
    10'd6:  neuron_4_mul_1_p <= Pix_34;
    10'd7:  neuron_4_mul_1_p <= Pix_35;
    10'd8:  neuron_4_mul_1_p <= Pix_36;
    10'd9:  neuron_4_mul_1_p <= Pix_37;
    10'd10:  neuron_4_mul_1_p <= Pix_38;
    10'd11:  neuron_4_mul_1_p <= Pix_39;
    10'd12:  neuron_4_mul_1_p <= Pix_40;
    10'd13:  neuron_4_mul_1_p <= Pix_41;
    10'd14:  neuron_4_mul_1_p <= Pix_42;
    10'd15:  neuron_4_mul_1_p <= Pix_43;
    10'd16:  neuron_4_mul_1_p <= Pix_44;
    10'd17:  neuron_4_mul_1_p <= Pix_45;
    10'd18:  neuron_4_mul_1_p <= Pix_46;
    10'd19:  neuron_4_mul_1_p <= Pix_47;
    10'd20:  neuron_4_mul_1_p <= Pix_48;
    10'd21:  neuron_4_mul_1_p <= Pix_49;
    10'd22:  neuron_4_mul_1_p <= Pix_50;
    10'd23:  neuron_4_mul_1_p <= Pix_51;
    10'd24:  neuron_4_mul_1_p <= Pix_52;
    10'd25:  neuron_4_mul_1_p <= Pix_53;
    10'd26:  neuron_4_mul_1_p <= Pix_54;
    10'd27:  neuron_4_mul_1_p <= Pix_55;
    default: neuron_4_mul_1_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_2_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_2_p <= Pix_56;
    10'd1:  neuron_4_mul_2_p <= Pix_57;
    10'd2:  neuron_4_mul_2_p <= Pix_58;
    10'd3:  neuron_4_mul_2_p <= Pix_59;
    10'd4:  neuron_4_mul_2_p <= Pix_60;
    10'd5:  neuron_4_mul_2_p <= Pix_61;
    10'd6:  neuron_4_mul_2_p <= Pix_62;
    10'd7:  neuron_4_mul_2_p <= Pix_63;
    10'd8:  neuron_4_mul_2_p <= Pix_64;
    10'd9:  neuron_4_mul_2_p <= Pix_65;
    10'd10:  neuron_4_mul_2_p <= Pix_66;
    10'd11:  neuron_4_mul_2_p <= Pix_67;
    10'd12:  neuron_4_mul_2_p <= Pix_68;
    10'd13:  neuron_4_mul_2_p <= Pix_69;
    10'd14:  neuron_4_mul_2_p <= Pix_70;
    10'd15:  neuron_4_mul_2_p <= Pix_71;
    10'd16:  neuron_4_mul_2_p <= Pix_72;
    10'd17:  neuron_4_mul_2_p <= Pix_73;
    10'd18:  neuron_4_mul_2_p <= Pix_74;
    10'd19:  neuron_4_mul_2_p <= Pix_75;
    10'd20:  neuron_4_mul_2_p <= Pix_76;
    10'd21:  neuron_4_mul_2_p <= Pix_77;
    10'd22:  neuron_4_mul_2_p <= Pix_78;
    10'd23:  neuron_4_mul_2_p <= Pix_79;
    10'd24:  neuron_4_mul_2_p <= Pix_80;
    10'd25:  neuron_4_mul_2_p <= Pix_81;
    10'd26:  neuron_4_mul_2_p <= Pix_82;
    10'd27:  neuron_4_mul_2_p <= Pix_83;
    default: neuron_4_mul_2_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_3_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_3_p <= Pix_84;
    10'd1:  neuron_4_mul_3_p <= Pix_85;
    10'd2:  neuron_4_mul_3_p <= Pix_86;
    10'd3:  neuron_4_mul_3_p <= Pix_87;
    10'd4:  neuron_4_mul_3_p <= Pix_88;
    10'd5:  neuron_4_mul_3_p <= Pix_89;
    10'd6:  neuron_4_mul_3_p <= Pix_90;
    10'd7:  neuron_4_mul_3_p <= Pix_91;
    10'd8:  neuron_4_mul_3_p <= Pix_92;
    10'd9:  neuron_4_mul_3_p <= Pix_93;
    10'd10:  neuron_4_mul_3_p <= Pix_94;
    10'd11:  neuron_4_mul_3_p <= Pix_95;
    10'd12:  neuron_4_mul_3_p <= Pix_96;
    10'd13:  neuron_4_mul_3_p <= Pix_97;
    10'd14:  neuron_4_mul_3_p <= Pix_98;
    10'd15:  neuron_4_mul_3_p <= Pix_99;
    10'd16:  neuron_4_mul_3_p <= Pix_100;
    10'd17:  neuron_4_mul_3_p <= Pix_101;
    10'd18:  neuron_4_mul_3_p <= Pix_102;
    10'd19:  neuron_4_mul_3_p <= Pix_103;
    10'd20:  neuron_4_mul_3_p <= Pix_104;
    10'd21:  neuron_4_mul_3_p <= Pix_105;
    10'd22:  neuron_4_mul_3_p <= Pix_106;
    10'd23:  neuron_4_mul_3_p <= Pix_107;
    10'd24:  neuron_4_mul_3_p <= Pix_108;
    10'd25:  neuron_4_mul_3_p <= Pix_109;
    10'd26:  neuron_4_mul_3_p <= Pix_110;
    10'd27:  neuron_4_mul_3_p <= Pix_111;
    default: neuron_4_mul_3_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_4_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_4_p <= Pix_112;
    10'd1:  neuron_4_mul_4_p <= Pix_113;
    10'd2:  neuron_4_mul_4_p <= Pix_114;
    10'd3:  neuron_4_mul_4_p <= Pix_115;
    10'd4:  neuron_4_mul_4_p <= Pix_116;
    10'd5:  neuron_4_mul_4_p <= Pix_117;
    10'd6:  neuron_4_mul_4_p <= Pix_118;
    10'd7:  neuron_4_mul_4_p <= Pix_119;
    10'd8:  neuron_4_mul_4_p <= Pix_120;
    10'd9:  neuron_4_mul_4_p <= Pix_121;
    10'd10:  neuron_4_mul_4_p <= Pix_122;
    10'd11:  neuron_4_mul_4_p <= Pix_123;
    10'd12:  neuron_4_mul_4_p <= Pix_124;
    10'd13:  neuron_4_mul_4_p <= Pix_125;
    10'd14:  neuron_4_mul_4_p <= Pix_126;
    10'd15:  neuron_4_mul_4_p <= Pix_127;
    10'd16:  neuron_4_mul_4_p <= Pix_128;
    10'd17:  neuron_4_mul_4_p <= Pix_129;
    10'd18:  neuron_4_mul_4_p <= Pix_130;
    10'd19:  neuron_4_mul_4_p <= Pix_131;
    10'd20:  neuron_4_mul_4_p <= Pix_132;
    10'd21:  neuron_4_mul_4_p <= Pix_133;
    10'd22:  neuron_4_mul_4_p <= Pix_134;
    10'd23:  neuron_4_mul_4_p <= Pix_135;
    10'd24:  neuron_4_mul_4_p <= Pix_136;
    10'd25:  neuron_4_mul_4_p <= Pix_137;
    10'd26:  neuron_4_mul_4_p <= Pix_138;
    10'd27:  neuron_4_mul_4_p <= Pix_139;
    default: neuron_4_mul_4_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_5_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_5_p <= Pix_140;
    10'd1:  neuron_4_mul_5_p <= Pix_141;
    10'd2:  neuron_4_mul_5_p <= Pix_142;
    10'd3:  neuron_4_mul_5_p <= Pix_143;
    10'd4:  neuron_4_mul_5_p <= Pix_144;
    10'd5:  neuron_4_mul_5_p <= Pix_145;
    10'd6:  neuron_4_mul_5_p <= Pix_146;
    10'd7:  neuron_4_mul_5_p <= Pix_147;
    10'd8:  neuron_4_mul_5_p <= Pix_148;
    10'd9:  neuron_4_mul_5_p <= Pix_149;
    10'd10:  neuron_4_mul_5_p <= Pix_150;
    10'd11:  neuron_4_mul_5_p <= Pix_151;
    10'd12:  neuron_4_mul_5_p <= Pix_152;
    10'd13:  neuron_4_mul_5_p <= Pix_153;
    10'd14:  neuron_4_mul_5_p <= Pix_154;
    10'd15:  neuron_4_mul_5_p <= Pix_155;
    10'd16:  neuron_4_mul_5_p <= Pix_156;
    10'd17:  neuron_4_mul_5_p <= Pix_157;
    10'd18:  neuron_4_mul_5_p <= Pix_158;
    10'd19:  neuron_4_mul_5_p <= Pix_159;
    10'd20:  neuron_4_mul_5_p <= Pix_160;
    10'd21:  neuron_4_mul_5_p <= Pix_161;
    10'd22:  neuron_4_mul_5_p <= Pix_162;
    10'd23:  neuron_4_mul_5_p <= Pix_163;
    10'd24:  neuron_4_mul_5_p <= Pix_164;
    10'd25:  neuron_4_mul_5_p <= Pix_165;
    10'd26:  neuron_4_mul_5_p <= Pix_166;
    10'd27:  neuron_4_mul_5_p <= Pix_167;
    default: neuron_4_mul_5_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_6_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_6_p <= Pix_168;
    10'd1:  neuron_4_mul_6_p <= Pix_169;
    10'd2:  neuron_4_mul_6_p <= Pix_170;
    10'd3:  neuron_4_mul_6_p <= Pix_171;
    10'd4:  neuron_4_mul_6_p <= Pix_172;
    10'd5:  neuron_4_mul_6_p <= Pix_173;
    10'd6:  neuron_4_mul_6_p <= Pix_174;
    10'd7:  neuron_4_mul_6_p <= Pix_175;
    10'd8:  neuron_4_mul_6_p <= Pix_176;
    10'd9:  neuron_4_mul_6_p <= Pix_177;
    10'd10:  neuron_4_mul_6_p <= Pix_178;
    10'd11:  neuron_4_mul_6_p <= Pix_179;
    10'd12:  neuron_4_mul_6_p <= Pix_180;
    10'd13:  neuron_4_mul_6_p <= Pix_181;
    10'd14:  neuron_4_mul_6_p <= Pix_182;
    10'd15:  neuron_4_mul_6_p <= Pix_183;
    10'd16:  neuron_4_mul_6_p <= Pix_184;
    10'd17:  neuron_4_mul_6_p <= Pix_185;
    10'd18:  neuron_4_mul_6_p <= Pix_186;
    10'd19:  neuron_4_mul_6_p <= Pix_187;
    10'd20:  neuron_4_mul_6_p <= Pix_188;
    10'd21:  neuron_4_mul_6_p <= Pix_189;
    10'd22:  neuron_4_mul_6_p <= Pix_190;
    10'd23:  neuron_4_mul_6_p <= Pix_191;
    10'd24:  neuron_4_mul_6_p <= Pix_192;
    10'd25:  neuron_4_mul_6_p <= Pix_193;
    10'd26:  neuron_4_mul_6_p <= Pix_194;
    10'd27:  neuron_4_mul_6_p <= Pix_195;
    default: neuron_4_mul_6_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_7_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_7_p <= Pix_196;
    10'd1:  neuron_4_mul_7_p <= Pix_197;
    10'd2:  neuron_4_mul_7_p <= Pix_198;
    10'd3:  neuron_4_mul_7_p <= Pix_199;
    10'd4:  neuron_4_mul_7_p <= Pix_200;
    10'd5:  neuron_4_mul_7_p <= Pix_201;
    10'd6:  neuron_4_mul_7_p <= Pix_202;
    10'd7:  neuron_4_mul_7_p <= Pix_203;
    10'd8:  neuron_4_mul_7_p <= Pix_204;
    10'd9:  neuron_4_mul_7_p <= Pix_205;
    10'd10:  neuron_4_mul_7_p <= Pix_206;
    10'd11:  neuron_4_mul_7_p <= Pix_207;
    10'd12:  neuron_4_mul_7_p <= Pix_208;
    10'd13:  neuron_4_mul_7_p <= Pix_209;
    10'd14:  neuron_4_mul_7_p <= Pix_210;
    10'd15:  neuron_4_mul_7_p <= Pix_211;
    10'd16:  neuron_4_mul_7_p <= Pix_212;
    10'd17:  neuron_4_mul_7_p <= Pix_213;
    10'd18:  neuron_4_mul_7_p <= Pix_214;
    10'd19:  neuron_4_mul_7_p <= Pix_215;
    10'd20:  neuron_4_mul_7_p <= Pix_216;
    10'd21:  neuron_4_mul_7_p <= Pix_217;
    10'd22:  neuron_4_mul_7_p <= Pix_218;
    10'd23:  neuron_4_mul_7_p <= Pix_219;
    10'd24:  neuron_4_mul_7_p <= Pix_220;
    10'd25:  neuron_4_mul_7_p <= Pix_221;
    10'd26:  neuron_4_mul_7_p <= Pix_222;
    10'd27:  neuron_4_mul_7_p <= Pix_223;
    default: neuron_4_mul_7_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_8_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_8_p <= Pix_224;
    10'd1:  neuron_4_mul_8_p <= Pix_225;
    10'd2:  neuron_4_mul_8_p <= Pix_226;
    10'd3:  neuron_4_mul_8_p <= Pix_227;
    10'd4:  neuron_4_mul_8_p <= Pix_228;
    10'd5:  neuron_4_mul_8_p <= Pix_229;
    10'd6:  neuron_4_mul_8_p <= Pix_230;
    10'd7:  neuron_4_mul_8_p <= Pix_231;
    10'd8:  neuron_4_mul_8_p <= Pix_232;
    10'd9:  neuron_4_mul_8_p <= Pix_233;
    10'd10:  neuron_4_mul_8_p <= Pix_234;
    10'd11:  neuron_4_mul_8_p <= Pix_235;
    10'd12:  neuron_4_mul_8_p <= Pix_236;
    10'd13:  neuron_4_mul_8_p <= Pix_237;
    10'd14:  neuron_4_mul_8_p <= Pix_238;
    10'd15:  neuron_4_mul_8_p <= Pix_239;
    10'd16:  neuron_4_mul_8_p <= Pix_240;
    10'd17:  neuron_4_mul_8_p <= Pix_241;
    10'd18:  neuron_4_mul_8_p <= Pix_242;
    10'd19:  neuron_4_mul_8_p <= Pix_243;
    10'd20:  neuron_4_mul_8_p <= Pix_244;
    10'd21:  neuron_4_mul_8_p <= Pix_245;
    10'd22:  neuron_4_mul_8_p <= Pix_246;
    10'd23:  neuron_4_mul_8_p <= Pix_247;
    10'd24:  neuron_4_mul_8_p <= Pix_248;
    10'd25:  neuron_4_mul_8_p <= Pix_249;
    10'd26:  neuron_4_mul_8_p <= Pix_250;
    10'd27:  neuron_4_mul_8_p <= Pix_251;
    default: neuron_4_mul_8_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_9_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_9_p <= Pix_252;
    10'd1:  neuron_4_mul_9_p <= Pix_253;
    10'd2:  neuron_4_mul_9_p <= Pix_254;
    10'd3:  neuron_4_mul_9_p <= Pix_255;
    10'd4:  neuron_4_mul_9_p <= Pix_256;
    10'd5:  neuron_4_mul_9_p <= Pix_257;
    10'd6:  neuron_4_mul_9_p <= Pix_258;
    10'd7:  neuron_4_mul_9_p <= Pix_259;
    10'd8:  neuron_4_mul_9_p <= Pix_260;
    10'd9:  neuron_4_mul_9_p <= Pix_261;
    10'd10:  neuron_4_mul_9_p <= Pix_262;
    10'd11:  neuron_4_mul_9_p <= Pix_263;
    10'd12:  neuron_4_mul_9_p <= Pix_264;
    10'd13:  neuron_4_mul_9_p <= Pix_265;
    10'd14:  neuron_4_mul_9_p <= Pix_266;
    10'd15:  neuron_4_mul_9_p <= Pix_267;
    10'd16:  neuron_4_mul_9_p <= Pix_268;
    10'd17:  neuron_4_mul_9_p <= Pix_269;
    10'd18:  neuron_4_mul_9_p <= Pix_270;
    10'd19:  neuron_4_mul_9_p <= Pix_271;
    10'd20:  neuron_4_mul_9_p <= Pix_272;
    10'd21:  neuron_4_mul_9_p <= Pix_273;
    10'd22:  neuron_4_mul_9_p <= Pix_274;
    10'd23:  neuron_4_mul_9_p <= Pix_275;
    10'd24:  neuron_4_mul_9_p <= Pix_276;
    10'd25:  neuron_4_mul_9_p <= Pix_277;
    10'd26:  neuron_4_mul_9_p <= Pix_278;
    10'd27:  neuron_4_mul_9_p <= Pix_279;
    default: neuron_4_mul_9_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_10_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_10_p <= Pix_280;
    10'd1:  neuron_4_mul_10_p <= Pix_281;
    10'd2:  neuron_4_mul_10_p <= Pix_282;
    10'd3:  neuron_4_mul_10_p <= Pix_283;
    10'd4:  neuron_4_mul_10_p <= Pix_284;
    10'd5:  neuron_4_mul_10_p <= Pix_285;
    10'd6:  neuron_4_mul_10_p <= Pix_286;
    10'd7:  neuron_4_mul_10_p <= Pix_287;
    10'd8:  neuron_4_mul_10_p <= Pix_288;
    10'd9:  neuron_4_mul_10_p <= Pix_289;
    10'd10:  neuron_4_mul_10_p <= Pix_290;
    10'd11:  neuron_4_mul_10_p <= Pix_291;
    10'd12:  neuron_4_mul_10_p <= Pix_292;
    10'd13:  neuron_4_mul_10_p <= Pix_293;
    10'd14:  neuron_4_mul_10_p <= Pix_294;
    10'd15:  neuron_4_mul_10_p <= Pix_295;
    10'd16:  neuron_4_mul_10_p <= Pix_296;
    10'd17:  neuron_4_mul_10_p <= Pix_297;
    10'd18:  neuron_4_mul_10_p <= Pix_298;
    10'd19:  neuron_4_mul_10_p <= Pix_299;
    10'd20:  neuron_4_mul_10_p <= Pix_300;
    10'd21:  neuron_4_mul_10_p <= Pix_301;
    10'd22:  neuron_4_mul_10_p <= Pix_302;
    10'd23:  neuron_4_mul_10_p <= Pix_303;
    10'd24:  neuron_4_mul_10_p <= Pix_304;
    10'd25:  neuron_4_mul_10_p <= Pix_305;
    10'd26:  neuron_4_mul_10_p <= Pix_306;
    10'd27:  neuron_4_mul_10_p <= Pix_307;
    default: neuron_4_mul_10_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_11_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_11_p <= Pix_308;
    10'd1:  neuron_4_mul_11_p <= Pix_309;
    10'd2:  neuron_4_mul_11_p <= Pix_310;
    10'd3:  neuron_4_mul_11_p <= Pix_311;
    10'd4:  neuron_4_mul_11_p <= Pix_312;
    10'd5:  neuron_4_mul_11_p <= Pix_313;
    10'd6:  neuron_4_mul_11_p <= Pix_314;
    10'd7:  neuron_4_mul_11_p <= Pix_315;
    10'd8:  neuron_4_mul_11_p <= Pix_316;
    10'd9:  neuron_4_mul_11_p <= Pix_317;
    10'd10:  neuron_4_mul_11_p <= Pix_318;
    10'd11:  neuron_4_mul_11_p <= Pix_319;
    10'd12:  neuron_4_mul_11_p <= Pix_320;
    10'd13:  neuron_4_mul_11_p <= Pix_321;
    10'd14:  neuron_4_mul_11_p <= Pix_322;
    10'd15:  neuron_4_mul_11_p <= Pix_323;
    10'd16:  neuron_4_mul_11_p <= Pix_324;
    10'd17:  neuron_4_mul_11_p <= Pix_325;
    10'd18:  neuron_4_mul_11_p <= Pix_326;
    10'd19:  neuron_4_mul_11_p <= Pix_327;
    10'd20:  neuron_4_mul_11_p <= Pix_328;
    10'd21:  neuron_4_mul_11_p <= Pix_329;
    10'd22:  neuron_4_mul_11_p <= Pix_330;
    10'd23:  neuron_4_mul_11_p <= Pix_331;
    10'd24:  neuron_4_mul_11_p <= Pix_332;
    10'd25:  neuron_4_mul_11_p <= Pix_333;
    10'd26:  neuron_4_mul_11_p <= Pix_334;
    10'd27:  neuron_4_mul_11_p <= Pix_335;
    default: neuron_4_mul_11_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_12_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_12_p <= Pix_336;
    10'd1:  neuron_4_mul_12_p <= Pix_337;
    10'd2:  neuron_4_mul_12_p <= Pix_338;
    10'd3:  neuron_4_mul_12_p <= Pix_339;
    10'd4:  neuron_4_mul_12_p <= Pix_340;
    10'd5:  neuron_4_mul_12_p <= Pix_341;
    10'd6:  neuron_4_mul_12_p <= Pix_342;
    10'd7:  neuron_4_mul_12_p <= Pix_343;
    10'd8:  neuron_4_mul_12_p <= Pix_344;
    10'd9:  neuron_4_mul_12_p <= Pix_345;
    10'd10:  neuron_4_mul_12_p <= Pix_346;
    10'd11:  neuron_4_mul_12_p <= Pix_347;
    10'd12:  neuron_4_mul_12_p <= Pix_348;
    10'd13:  neuron_4_mul_12_p <= Pix_349;
    10'd14:  neuron_4_mul_12_p <= Pix_350;
    10'd15:  neuron_4_mul_12_p <= Pix_351;
    10'd16:  neuron_4_mul_12_p <= Pix_352;
    10'd17:  neuron_4_mul_12_p <= Pix_353;
    10'd18:  neuron_4_mul_12_p <= Pix_354;
    10'd19:  neuron_4_mul_12_p <= Pix_355;
    10'd20:  neuron_4_mul_12_p <= Pix_356;
    10'd21:  neuron_4_mul_12_p <= Pix_357;
    10'd22:  neuron_4_mul_12_p <= Pix_358;
    10'd23:  neuron_4_mul_12_p <= Pix_359;
    10'd24:  neuron_4_mul_12_p <= Pix_360;
    10'd25:  neuron_4_mul_12_p <= Pix_361;
    10'd26:  neuron_4_mul_12_p <= Pix_362;
    10'd27:  neuron_4_mul_12_p <= Pix_363;
    default: neuron_4_mul_12_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_13_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_13_p <= Pix_364;
    10'd1:  neuron_4_mul_13_p <= Pix_365;
    10'd2:  neuron_4_mul_13_p <= Pix_366;
    10'd3:  neuron_4_mul_13_p <= Pix_367;
    10'd4:  neuron_4_mul_13_p <= Pix_368;
    10'd5:  neuron_4_mul_13_p <= Pix_369;
    10'd6:  neuron_4_mul_13_p <= Pix_370;
    10'd7:  neuron_4_mul_13_p <= Pix_371;
    10'd8:  neuron_4_mul_13_p <= Pix_372;
    10'd9:  neuron_4_mul_13_p <= Pix_373;
    10'd10:  neuron_4_mul_13_p <= Pix_374;
    10'd11:  neuron_4_mul_13_p <= Pix_375;
    10'd12:  neuron_4_mul_13_p <= Pix_376;
    10'd13:  neuron_4_mul_13_p <= Pix_377;
    10'd14:  neuron_4_mul_13_p <= Pix_378;
    10'd15:  neuron_4_mul_13_p <= Pix_379;
    10'd16:  neuron_4_mul_13_p <= Pix_380;
    10'd17:  neuron_4_mul_13_p <= Pix_381;
    10'd18:  neuron_4_mul_13_p <= Pix_382;
    10'd19:  neuron_4_mul_13_p <= Pix_383;
    10'd20:  neuron_4_mul_13_p <= Pix_384;
    10'd21:  neuron_4_mul_13_p <= Pix_385;
    10'd22:  neuron_4_mul_13_p <= Pix_386;
    10'd23:  neuron_4_mul_13_p <= Pix_387;
    10'd24:  neuron_4_mul_13_p <= Pix_388;
    10'd25:  neuron_4_mul_13_p <= Pix_389;
    10'd26:  neuron_4_mul_13_p <= Pix_390;
    10'd27:  neuron_4_mul_13_p <= Pix_391;
    default: neuron_4_mul_13_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_14_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_14_p <= Pix_392;
    10'd1:  neuron_4_mul_14_p <= Pix_393;
    10'd2:  neuron_4_mul_14_p <= Pix_394;
    10'd3:  neuron_4_mul_14_p <= Pix_395;
    10'd4:  neuron_4_mul_14_p <= Pix_396;
    10'd5:  neuron_4_mul_14_p <= Pix_397;
    10'd6:  neuron_4_mul_14_p <= Pix_398;
    10'd7:  neuron_4_mul_14_p <= Pix_399;
    10'd8:  neuron_4_mul_14_p <= Pix_400;
    10'd9:  neuron_4_mul_14_p <= Pix_401;
    10'd10:  neuron_4_mul_14_p <= Pix_402;
    10'd11:  neuron_4_mul_14_p <= Pix_403;
    10'd12:  neuron_4_mul_14_p <= Pix_404;
    10'd13:  neuron_4_mul_14_p <= Pix_405;
    10'd14:  neuron_4_mul_14_p <= Pix_406;
    10'd15:  neuron_4_mul_14_p <= Pix_407;
    10'd16:  neuron_4_mul_14_p <= Pix_408;
    10'd17:  neuron_4_mul_14_p <= Pix_409;
    10'd18:  neuron_4_mul_14_p <= Pix_410;
    10'd19:  neuron_4_mul_14_p <= Pix_411;
    10'd20:  neuron_4_mul_14_p <= Pix_412;
    10'd21:  neuron_4_mul_14_p <= Pix_413;
    10'd22:  neuron_4_mul_14_p <= Pix_414;
    10'd23:  neuron_4_mul_14_p <= Pix_415;
    10'd24:  neuron_4_mul_14_p <= Pix_416;
    10'd25:  neuron_4_mul_14_p <= Pix_417;
    10'd26:  neuron_4_mul_14_p <= Pix_418;
    10'd27:  neuron_4_mul_14_p <= Pix_419;
    default: neuron_4_mul_14_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_15_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_15_p <= Pix_420;
    10'd1:  neuron_4_mul_15_p <= Pix_421;
    10'd2:  neuron_4_mul_15_p <= Pix_422;
    10'd3:  neuron_4_mul_15_p <= Pix_423;
    10'd4:  neuron_4_mul_15_p <= Pix_424;
    10'd5:  neuron_4_mul_15_p <= Pix_425;
    10'd6:  neuron_4_mul_15_p <= Pix_426;
    10'd7:  neuron_4_mul_15_p <= Pix_427;
    10'd8:  neuron_4_mul_15_p <= Pix_428;
    10'd9:  neuron_4_mul_15_p <= Pix_429;
    10'd10:  neuron_4_mul_15_p <= Pix_430;
    10'd11:  neuron_4_mul_15_p <= Pix_431;
    10'd12:  neuron_4_mul_15_p <= Pix_432;
    10'd13:  neuron_4_mul_15_p <= Pix_433;
    10'd14:  neuron_4_mul_15_p <= Pix_434;
    10'd15:  neuron_4_mul_15_p <= Pix_435;
    10'd16:  neuron_4_mul_15_p <= Pix_436;
    10'd17:  neuron_4_mul_15_p <= Pix_437;
    10'd18:  neuron_4_mul_15_p <= Pix_438;
    10'd19:  neuron_4_mul_15_p <= Pix_439;
    10'd20:  neuron_4_mul_15_p <= Pix_440;
    10'd21:  neuron_4_mul_15_p <= Pix_441;
    10'd22:  neuron_4_mul_15_p <= Pix_442;
    10'd23:  neuron_4_mul_15_p <= Pix_443;
    10'd24:  neuron_4_mul_15_p <= Pix_444;
    10'd25:  neuron_4_mul_15_p <= Pix_445;
    10'd26:  neuron_4_mul_15_p <= Pix_446;
    10'd27:  neuron_4_mul_15_p <= Pix_447;
    default: neuron_4_mul_15_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_16_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_16_p <= Pix_448;
    10'd1:  neuron_4_mul_16_p <= Pix_449;
    10'd2:  neuron_4_mul_16_p <= Pix_450;
    10'd3:  neuron_4_mul_16_p <= Pix_451;
    10'd4:  neuron_4_mul_16_p <= Pix_452;
    10'd5:  neuron_4_mul_16_p <= Pix_453;
    10'd6:  neuron_4_mul_16_p <= Pix_454;
    10'd7:  neuron_4_mul_16_p <= Pix_455;
    10'd8:  neuron_4_mul_16_p <= Pix_456;
    10'd9:  neuron_4_mul_16_p <= Pix_457;
    10'd10:  neuron_4_mul_16_p <= Pix_458;
    10'd11:  neuron_4_mul_16_p <= Pix_459;
    10'd12:  neuron_4_mul_16_p <= Pix_460;
    10'd13:  neuron_4_mul_16_p <= Pix_461;
    10'd14:  neuron_4_mul_16_p <= Pix_462;
    10'd15:  neuron_4_mul_16_p <= Pix_463;
    10'd16:  neuron_4_mul_16_p <= Pix_464;
    10'd17:  neuron_4_mul_16_p <= Pix_465;
    10'd18:  neuron_4_mul_16_p <= Pix_466;
    10'd19:  neuron_4_mul_16_p <= Pix_467;
    10'd20:  neuron_4_mul_16_p <= Pix_468;
    10'd21:  neuron_4_mul_16_p <= Pix_469;
    10'd22:  neuron_4_mul_16_p <= Pix_470;
    10'd23:  neuron_4_mul_16_p <= Pix_471;
    10'd24:  neuron_4_mul_16_p <= Pix_472;
    10'd25:  neuron_4_mul_16_p <= Pix_473;
    10'd26:  neuron_4_mul_16_p <= Pix_474;
    10'd27:  neuron_4_mul_16_p <= Pix_475;
    default: neuron_4_mul_16_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_17_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_17_p <= Pix_476;
    10'd1:  neuron_4_mul_17_p <= Pix_477;
    10'd2:  neuron_4_mul_17_p <= Pix_478;
    10'd3:  neuron_4_mul_17_p <= Pix_479;
    10'd4:  neuron_4_mul_17_p <= Pix_480;
    10'd5:  neuron_4_mul_17_p <= Pix_481;
    10'd6:  neuron_4_mul_17_p <= Pix_482;
    10'd7:  neuron_4_mul_17_p <= Pix_483;
    10'd8:  neuron_4_mul_17_p <= Pix_484;
    10'd9:  neuron_4_mul_17_p <= Pix_485;
    10'd10:  neuron_4_mul_17_p <= Pix_486;
    10'd11:  neuron_4_mul_17_p <= Pix_487;
    10'd12:  neuron_4_mul_17_p <= Pix_488;
    10'd13:  neuron_4_mul_17_p <= Pix_489;
    10'd14:  neuron_4_mul_17_p <= Pix_490;
    10'd15:  neuron_4_mul_17_p <= Pix_491;
    10'd16:  neuron_4_mul_17_p <= Pix_492;
    10'd17:  neuron_4_mul_17_p <= Pix_493;
    10'd18:  neuron_4_mul_17_p <= Pix_494;
    10'd19:  neuron_4_mul_17_p <= Pix_495;
    10'd20:  neuron_4_mul_17_p <= Pix_496;
    10'd21:  neuron_4_mul_17_p <= Pix_497;
    10'd22:  neuron_4_mul_17_p <= Pix_498;
    10'd23:  neuron_4_mul_17_p <= Pix_499;
    10'd24:  neuron_4_mul_17_p <= Pix_500;
    10'd25:  neuron_4_mul_17_p <= Pix_501;
    10'd26:  neuron_4_mul_17_p <= Pix_502;
    10'd27:  neuron_4_mul_17_p <= Pix_503;
    default: neuron_4_mul_17_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_18_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_18_p <= Pix_504;
    10'd1:  neuron_4_mul_18_p <= Pix_505;
    10'd2:  neuron_4_mul_18_p <= Pix_506;
    10'd3:  neuron_4_mul_18_p <= Pix_507;
    10'd4:  neuron_4_mul_18_p <= Pix_508;
    10'd5:  neuron_4_mul_18_p <= Pix_509;
    10'd6:  neuron_4_mul_18_p <= Pix_510;
    10'd7:  neuron_4_mul_18_p <= Pix_511;
    10'd8:  neuron_4_mul_18_p <= Pix_512;
    10'd9:  neuron_4_mul_18_p <= Pix_513;
    10'd10:  neuron_4_mul_18_p <= Pix_514;
    10'd11:  neuron_4_mul_18_p <= Pix_515;
    10'd12:  neuron_4_mul_18_p <= Pix_516;
    10'd13:  neuron_4_mul_18_p <= Pix_517;
    10'd14:  neuron_4_mul_18_p <= Pix_518;
    10'd15:  neuron_4_mul_18_p <= Pix_519;
    10'd16:  neuron_4_mul_18_p <= Pix_520;
    10'd17:  neuron_4_mul_18_p <= Pix_521;
    10'd18:  neuron_4_mul_18_p <= Pix_522;
    10'd19:  neuron_4_mul_18_p <= Pix_523;
    10'd20:  neuron_4_mul_18_p <= Pix_524;
    10'd21:  neuron_4_mul_18_p <= Pix_525;
    10'd22:  neuron_4_mul_18_p <= Pix_526;
    10'd23:  neuron_4_mul_18_p <= Pix_527;
    10'd24:  neuron_4_mul_18_p <= Pix_528;
    10'd25:  neuron_4_mul_18_p <= Pix_529;
    10'd26:  neuron_4_mul_18_p <= Pix_530;
    10'd27:  neuron_4_mul_18_p <= Pix_531;
    default: neuron_4_mul_18_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_19_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_19_p <= Pix_532;
    10'd1:  neuron_4_mul_19_p <= Pix_533;
    10'd2:  neuron_4_mul_19_p <= Pix_534;
    10'd3:  neuron_4_mul_19_p <= Pix_535;
    10'd4:  neuron_4_mul_19_p <= Pix_536;
    10'd5:  neuron_4_mul_19_p <= Pix_537;
    10'd6:  neuron_4_mul_19_p <= Pix_538;
    10'd7:  neuron_4_mul_19_p <= Pix_539;
    10'd8:  neuron_4_mul_19_p <= Pix_540;
    10'd9:  neuron_4_mul_19_p <= Pix_541;
    10'd10:  neuron_4_mul_19_p <= Pix_542;
    10'd11:  neuron_4_mul_19_p <= Pix_543;
    10'd12:  neuron_4_mul_19_p <= Pix_544;
    10'd13:  neuron_4_mul_19_p <= Pix_545;
    10'd14:  neuron_4_mul_19_p <= Pix_546;
    10'd15:  neuron_4_mul_19_p <= Pix_547;
    10'd16:  neuron_4_mul_19_p <= Pix_548;
    10'd17:  neuron_4_mul_19_p <= Pix_549;
    10'd18:  neuron_4_mul_19_p <= Pix_550;
    10'd19:  neuron_4_mul_19_p <= Pix_551;
    10'd20:  neuron_4_mul_19_p <= Pix_552;
    10'd21:  neuron_4_mul_19_p <= Pix_553;
    10'd22:  neuron_4_mul_19_p <= Pix_554;
    10'd23:  neuron_4_mul_19_p <= Pix_555;
    10'd24:  neuron_4_mul_19_p <= Pix_556;
    10'd25:  neuron_4_mul_19_p <= Pix_557;
    10'd26:  neuron_4_mul_19_p <= Pix_558;
    10'd27:  neuron_4_mul_19_p <= Pix_559;
    default: neuron_4_mul_19_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_20_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_20_p <= Pix_560;
    10'd1:  neuron_4_mul_20_p <= Pix_561;
    10'd2:  neuron_4_mul_20_p <= Pix_562;
    10'd3:  neuron_4_mul_20_p <= Pix_563;
    10'd4:  neuron_4_mul_20_p <= Pix_564;
    10'd5:  neuron_4_mul_20_p <= Pix_565;
    10'd6:  neuron_4_mul_20_p <= Pix_566;
    10'd7:  neuron_4_mul_20_p <= Pix_567;
    10'd8:  neuron_4_mul_20_p <= Pix_568;
    10'd9:  neuron_4_mul_20_p <= Pix_569;
    10'd10:  neuron_4_mul_20_p <= Pix_570;
    10'd11:  neuron_4_mul_20_p <= Pix_571;
    10'd12:  neuron_4_mul_20_p <= Pix_572;
    10'd13:  neuron_4_mul_20_p <= Pix_573;
    10'd14:  neuron_4_mul_20_p <= Pix_574;
    10'd15:  neuron_4_mul_20_p <= Pix_575;
    10'd16:  neuron_4_mul_20_p <= Pix_576;
    10'd17:  neuron_4_mul_20_p <= Pix_577;
    10'd18:  neuron_4_mul_20_p <= Pix_578;
    10'd19:  neuron_4_mul_20_p <= Pix_579;
    10'd20:  neuron_4_mul_20_p <= Pix_580;
    10'd21:  neuron_4_mul_20_p <= Pix_581;
    10'd22:  neuron_4_mul_20_p <= Pix_582;
    10'd23:  neuron_4_mul_20_p <= Pix_583;
    10'd24:  neuron_4_mul_20_p <= Pix_584;
    10'd25:  neuron_4_mul_20_p <= Pix_585;
    10'd26:  neuron_4_mul_20_p <= Pix_586;
    10'd27:  neuron_4_mul_20_p <= Pix_587;
    default: neuron_4_mul_20_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_21_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_21_p <= Pix_588;
    10'd1:  neuron_4_mul_21_p <= Pix_589;
    10'd2:  neuron_4_mul_21_p <= Pix_590;
    10'd3:  neuron_4_mul_21_p <= Pix_591;
    10'd4:  neuron_4_mul_21_p <= Pix_592;
    10'd5:  neuron_4_mul_21_p <= Pix_593;
    10'd6:  neuron_4_mul_21_p <= Pix_594;
    10'd7:  neuron_4_mul_21_p <= Pix_595;
    10'd8:  neuron_4_mul_21_p <= Pix_596;
    10'd9:  neuron_4_mul_21_p <= Pix_597;
    10'd10:  neuron_4_mul_21_p <= Pix_598;
    10'd11:  neuron_4_mul_21_p <= Pix_599;
    10'd12:  neuron_4_mul_21_p <= Pix_600;
    10'd13:  neuron_4_mul_21_p <= Pix_601;
    10'd14:  neuron_4_mul_21_p <= Pix_602;
    10'd15:  neuron_4_mul_21_p <= Pix_603;
    10'd16:  neuron_4_mul_21_p <= Pix_604;
    10'd17:  neuron_4_mul_21_p <= Pix_605;
    10'd18:  neuron_4_mul_21_p <= Pix_606;
    10'd19:  neuron_4_mul_21_p <= Pix_607;
    10'd20:  neuron_4_mul_21_p <= Pix_608;
    10'd21:  neuron_4_mul_21_p <= Pix_609;
    10'd22:  neuron_4_mul_21_p <= Pix_610;
    10'd23:  neuron_4_mul_21_p <= Pix_611;
    10'd24:  neuron_4_mul_21_p <= Pix_612;
    10'd25:  neuron_4_mul_21_p <= Pix_613;
    10'd26:  neuron_4_mul_21_p <= Pix_614;
    10'd27:  neuron_4_mul_21_p <= Pix_615;
    default: neuron_4_mul_21_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_22_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_22_p <= Pix_616;
    10'd1:  neuron_4_mul_22_p <= Pix_617;
    10'd2:  neuron_4_mul_22_p <= Pix_618;
    10'd3:  neuron_4_mul_22_p <= Pix_619;
    10'd4:  neuron_4_mul_22_p <= Pix_620;
    10'd5:  neuron_4_mul_22_p <= Pix_621;
    10'd6:  neuron_4_mul_22_p <= Pix_622;
    10'd7:  neuron_4_mul_22_p <= Pix_623;
    10'd8:  neuron_4_mul_22_p <= Pix_624;
    10'd9:  neuron_4_mul_22_p <= Pix_625;
    10'd10:  neuron_4_mul_22_p <= Pix_626;
    10'd11:  neuron_4_mul_22_p <= Pix_627;
    10'd12:  neuron_4_mul_22_p <= Pix_628;
    10'd13:  neuron_4_mul_22_p <= Pix_629;
    10'd14:  neuron_4_mul_22_p <= Pix_630;
    10'd15:  neuron_4_mul_22_p <= Pix_631;
    10'd16:  neuron_4_mul_22_p <= Pix_632;
    10'd17:  neuron_4_mul_22_p <= Pix_633;
    10'd18:  neuron_4_mul_22_p <= Pix_634;
    10'd19:  neuron_4_mul_22_p <= Pix_635;
    10'd20:  neuron_4_mul_22_p <= Pix_636;
    10'd21:  neuron_4_mul_22_p <= Pix_637;
    10'd22:  neuron_4_mul_22_p <= Pix_638;
    10'd23:  neuron_4_mul_22_p <= Pix_639;
    10'd24:  neuron_4_mul_22_p <= Pix_640;
    10'd25:  neuron_4_mul_22_p <= Pix_641;
    10'd26:  neuron_4_mul_22_p <= Pix_642;
    10'd27:  neuron_4_mul_22_p <= Pix_643;
    default: neuron_4_mul_22_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_23_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_23_p <= Pix_644;
    10'd1:  neuron_4_mul_23_p <= Pix_645;
    10'd2:  neuron_4_mul_23_p <= Pix_646;
    10'd3:  neuron_4_mul_23_p <= Pix_647;
    10'd4:  neuron_4_mul_23_p <= Pix_648;
    10'd5:  neuron_4_mul_23_p <= Pix_649;
    10'd6:  neuron_4_mul_23_p <= Pix_650;
    10'd7:  neuron_4_mul_23_p <= Pix_651;
    10'd8:  neuron_4_mul_23_p <= Pix_652;
    10'd9:  neuron_4_mul_23_p <= Pix_653;
    10'd10:  neuron_4_mul_23_p <= Pix_654;
    10'd11:  neuron_4_mul_23_p <= Pix_655;
    10'd12:  neuron_4_mul_23_p <= Pix_656;
    10'd13:  neuron_4_mul_23_p <= Pix_657;
    10'd14:  neuron_4_mul_23_p <= Pix_658;
    10'd15:  neuron_4_mul_23_p <= Pix_659;
    10'd16:  neuron_4_mul_23_p <= Pix_660;
    10'd17:  neuron_4_mul_23_p <= Pix_661;
    10'd18:  neuron_4_mul_23_p <= Pix_662;
    10'd19:  neuron_4_mul_23_p <= Pix_663;
    10'd20:  neuron_4_mul_23_p <= Pix_664;
    10'd21:  neuron_4_mul_23_p <= Pix_665;
    10'd22:  neuron_4_mul_23_p <= Pix_666;
    10'd23:  neuron_4_mul_23_p <= Pix_667;
    10'd24:  neuron_4_mul_23_p <= Pix_668;
    10'd25:  neuron_4_mul_23_p <= Pix_669;
    10'd26:  neuron_4_mul_23_p <= Pix_670;
    10'd27:  neuron_4_mul_23_p <= Pix_671;
    default: neuron_4_mul_23_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_24_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_24_p <= Pix_672;
    10'd1:  neuron_4_mul_24_p <= Pix_673;
    10'd2:  neuron_4_mul_24_p <= Pix_674;
    10'd3:  neuron_4_mul_24_p <= Pix_675;
    10'd4:  neuron_4_mul_24_p <= Pix_676;
    10'd5:  neuron_4_mul_24_p <= Pix_677;
    10'd6:  neuron_4_mul_24_p <= Pix_678;
    10'd7:  neuron_4_mul_24_p <= Pix_679;
    10'd8:  neuron_4_mul_24_p <= Pix_680;
    10'd9:  neuron_4_mul_24_p <= Pix_681;
    10'd10:  neuron_4_mul_24_p <= Pix_682;
    10'd11:  neuron_4_mul_24_p <= Pix_683;
    10'd12:  neuron_4_mul_24_p <= Pix_684;
    10'd13:  neuron_4_mul_24_p <= Pix_685;
    10'd14:  neuron_4_mul_24_p <= Pix_686;
    10'd15:  neuron_4_mul_24_p <= Pix_687;
    10'd16:  neuron_4_mul_24_p <= Pix_688;
    10'd17:  neuron_4_mul_24_p <= Pix_689;
    10'd18:  neuron_4_mul_24_p <= Pix_690;
    10'd19:  neuron_4_mul_24_p <= Pix_691;
    10'd20:  neuron_4_mul_24_p <= Pix_692;
    10'd21:  neuron_4_mul_24_p <= Pix_693;
    10'd22:  neuron_4_mul_24_p <= Pix_694;
    10'd23:  neuron_4_mul_24_p <= Pix_695;
    10'd24:  neuron_4_mul_24_p <= Pix_696;
    10'd25:  neuron_4_mul_24_p <= Pix_697;
    10'd26:  neuron_4_mul_24_p <= Pix_698;
    10'd27:  neuron_4_mul_24_p <= Pix_699;
    default: neuron_4_mul_24_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_25_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_25_p <= Pix_700;
    10'd1:  neuron_4_mul_25_p <= Pix_701;
    10'd2:  neuron_4_mul_25_p <= Pix_702;
    10'd3:  neuron_4_mul_25_p <= Pix_703;
    10'd4:  neuron_4_mul_25_p <= Pix_704;
    10'd5:  neuron_4_mul_25_p <= Pix_705;
    10'd6:  neuron_4_mul_25_p <= Pix_706;
    10'd7:  neuron_4_mul_25_p <= Pix_707;
    10'd8:  neuron_4_mul_25_p <= Pix_708;
    10'd9:  neuron_4_mul_25_p <= Pix_709;
    10'd10:  neuron_4_mul_25_p <= Pix_710;
    10'd11:  neuron_4_mul_25_p <= Pix_711;
    10'd12:  neuron_4_mul_25_p <= Pix_712;
    10'd13:  neuron_4_mul_25_p <= Pix_713;
    10'd14:  neuron_4_mul_25_p <= Pix_714;
    10'd15:  neuron_4_mul_25_p <= Pix_715;
    10'd16:  neuron_4_mul_25_p <= Pix_716;
    10'd17:  neuron_4_mul_25_p <= Pix_717;
    10'd18:  neuron_4_mul_25_p <= Pix_718;
    10'd19:  neuron_4_mul_25_p <= Pix_719;
    10'd20:  neuron_4_mul_25_p <= Pix_720;
    10'd21:  neuron_4_mul_25_p <= Pix_721;
    10'd22:  neuron_4_mul_25_p <= Pix_722;
    10'd23:  neuron_4_mul_25_p <= Pix_723;
    10'd24:  neuron_4_mul_25_p <= Pix_724;
    10'd25:  neuron_4_mul_25_p <= Pix_725;
    10'd26:  neuron_4_mul_25_p <= Pix_726;
    10'd27:  neuron_4_mul_25_p <= Pix_727;
    default: neuron_4_mul_25_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_26_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_26_p <= Pix_728;
    10'd1:  neuron_4_mul_26_p <= Pix_729;
    10'd2:  neuron_4_mul_26_p <= Pix_730;
    10'd3:  neuron_4_mul_26_p <= Pix_731;
    10'd4:  neuron_4_mul_26_p <= Pix_732;
    10'd5:  neuron_4_mul_26_p <= Pix_733;
    10'd6:  neuron_4_mul_26_p <= Pix_734;
    10'd7:  neuron_4_mul_26_p <= Pix_735;
    10'd8:  neuron_4_mul_26_p <= Pix_736;
    10'd9:  neuron_4_mul_26_p <= Pix_737;
    10'd10:  neuron_4_mul_26_p <= Pix_738;
    10'd11:  neuron_4_mul_26_p <= Pix_739;
    10'd12:  neuron_4_mul_26_p <= Pix_740;
    10'd13:  neuron_4_mul_26_p <= Pix_741;
    10'd14:  neuron_4_mul_26_p <= Pix_742;
    10'd15:  neuron_4_mul_26_p <= Pix_743;
    10'd16:  neuron_4_mul_26_p <= Pix_744;
    10'd17:  neuron_4_mul_26_p <= Pix_745;
    10'd18:  neuron_4_mul_26_p <= Pix_746;
    10'd19:  neuron_4_mul_26_p <= Pix_747;
    10'd20:  neuron_4_mul_26_p <= Pix_748;
    10'd21:  neuron_4_mul_26_p <= Pix_749;
    10'd22:  neuron_4_mul_26_p <= Pix_750;
    10'd23:  neuron_4_mul_26_p <= Pix_751;
    10'd24:  neuron_4_mul_26_p <= Pix_752;
    10'd25:  neuron_4_mul_26_p <= Pix_753;
    10'd26:  neuron_4_mul_26_p <= Pix_754;
    10'd27:  neuron_4_mul_26_p <= Pix_755;
    default: neuron_4_mul_26_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_4_mul_27_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_4_mul_27_p <= Pix_756;
    10'd1:  neuron_4_mul_27_p <= Pix_757;
    10'd2:  neuron_4_mul_27_p <= Pix_758;
    10'd3:  neuron_4_mul_27_p <= Pix_759;
    10'd4:  neuron_4_mul_27_p <= Pix_760;
    10'd5:  neuron_4_mul_27_p <= Pix_761;
    10'd6:  neuron_4_mul_27_p <= Pix_762;
    10'd7:  neuron_4_mul_27_p <= Pix_763;
    10'd8:  neuron_4_mul_27_p <= Pix_764;
    10'd9:  neuron_4_mul_27_p <= Pix_765;
    10'd10:  neuron_4_mul_27_p <= Pix_766;
    10'd11:  neuron_4_mul_27_p <= Pix_767;
    10'd12:  neuron_4_mul_27_p <= Pix_768;
    10'd13:  neuron_4_mul_27_p <= Pix_769;
    10'd14:  neuron_4_mul_27_p <= Pix_770;
    10'd15:  neuron_4_mul_27_p <= Pix_771;
    10'd16:  neuron_4_mul_27_p <= Pix_772;
    10'd17:  neuron_4_mul_27_p <= Pix_773;
    10'd18:  neuron_4_mul_27_p <= Pix_774;
    10'd19:  neuron_4_mul_27_p <= Pix_775;
    10'd20:  neuron_4_mul_27_p <= Pix_776;
    10'd21:  neuron_4_mul_27_p <= Pix_777;
    10'd22:  neuron_4_mul_27_p <= Pix_778;
    10'd23:  neuron_4_mul_27_p <= Pix_779;
    10'd24:  neuron_4_mul_27_p <= Pix_780;
    10'd25:  neuron_4_mul_27_p <= Pix_781;
    10'd26:  neuron_4_mul_27_p <= Pix_782;
    10'd27:  neuron_4_mul_27_p <= Pix_783;
    default: neuron_4_mul_27_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_0_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_0_p <= Pix_0;
    10'd1:  neuron_5_mul_0_p <= Pix_1;
    10'd2:  neuron_5_mul_0_p <= Pix_2;
    10'd3:  neuron_5_mul_0_p <= Pix_3;
    10'd4:  neuron_5_mul_0_p <= Pix_4;
    10'd5:  neuron_5_mul_0_p <= Pix_5;
    10'd6:  neuron_5_mul_0_p <= Pix_6;
    10'd7:  neuron_5_mul_0_p <= Pix_7;
    10'd8:  neuron_5_mul_0_p <= Pix_8;
    10'd9:  neuron_5_mul_0_p <= Pix_9;
    10'd10:  neuron_5_mul_0_p <= Pix_10;
    10'd11:  neuron_5_mul_0_p <= Pix_11;
    10'd12:  neuron_5_mul_0_p <= Pix_12;
    10'd13:  neuron_5_mul_0_p <= Pix_13;
    10'd14:  neuron_5_mul_0_p <= Pix_14;
    10'd15:  neuron_5_mul_0_p <= Pix_15;
    10'd16:  neuron_5_mul_0_p <= Pix_16;
    10'd17:  neuron_5_mul_0_p <= Pix_17;
    10'd18:  neuron_5_mul_0_p <= Pix_18;
    10'd19:  neuron_5_mul_0_p <= Pix_19;
    10'd20:  neuron_5_mul_0_p <= Pix_20;
    10'd21:  neuron_5_mul_0_p <= Pix_21;
    10'd22:  neuron_5_mul_0_p <= Pix_22;
    10'd23:  neuron_5_mul_0_p <= Pix_23;
    10'd24:  neuron_5_mul_0_p <= Pix_24;
    10'd25:  neuron_5_mul_0_p <= Pix_25;
    10'd26:  neuron_5_mul_0_p <= Pix_26;
    10'd27:  neuron_5_mul_0_p <= Pix_27;
    default: neuron_5_mul_0_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_1_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_1_p <= Pix_28;
    10'd1:  neuron_5_mul_1_p <= Pix_29;
    10'd2:  neuron_5_mul_1_p <= Pix_30;
    10'd3:  neuron_5_mul_1_p <= Pix_31;
    10'd4:  neuron_5_mul_1_p <= Pix_32;
    10'd5:  neuron_5_mul_1_p <= Pix_33;
    10'd6:  neuron_5_mul_1_p <= Pix_34;
    10'd7:  neuron_5_mul_1_p <= Pix_35;
    10'd8:  neuron_5_mul_1_p <= Pix_36;
    10'd9:  neuron_5_mul_1_p <= Pix_37;
    10'd10:  neuron_5_mul_1_p <= Pix_38;
    10'd11:  neuron_5_mul_1_p <= Pix_39;
    10'd12:  neuron_5_mul_1_p <= Pix_40;
    10'd13:  neuron_5_mul_1_p <= Pix_41;
    10'd14:  neuron_5_mul_1_p <= Pix_42;
    10'd15:  neuron_5_mul_1_p <= Pix_43;
    10'd16:  neuron_5_mul_1_p <= Pix_44;
    10'd17:  neuron_5_mul_1_p <= Pix_45;
    10'd18:  neuron_5_mul_1_p <= Pix_46;
    10'd19:  neuron_5_mul_1_p <= Pix_47;
    10'd20:  neuron_5_mul_1_p <= Pix_48;
    10'd21:  neuron_5_mul_1_p <= Pix_49;
    10'd22:  neuron_5_mul_1_p <= Pix_50;
    10'd23:  neuron_5_mul_1_p <= Pix_51;
    10'd24:  neuron_5_mul_1_p <= Pix_52;
    10'd25:  neuron_5_mul_1_p <= Pix_53;
    10'd26:  neuron_5_mul_1_p <= Pix_54;
    10'd27:  neuron_5_mul_1_p <= Pix_55;
    default: neuron_5_mul_1_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_2_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_2_p <= Pix_56;
    10'd1:  neuron_5_mul_2_p <= Pix_57;
    10'd2:  neuron_5_mul_2_p <= Pix_58;
    10'd3:  neuron_5_mul_2_p <= Pix_59;
    10'd4:  neuron_5_mul_2_p <= Pix_60;
    10'd5:  neuron_5_mul_2_p <= Pix_61;
    10'd6:  neuron_5_mul_2_p <= Pix_62;
    10'd7:  neuron_5_mul_2_p <= Pix_63;
    10'd8:  neuron_5_mul_2_p <= Pix_64;
    10'd9:  neuron_5_mul_2_p <= Pix_65;
    10'd10:  neuron_5_mul_2_p <= Pix_66;
    10'd11:  neuron_5_mul_2_p <= Pix_67;
    10'd12:  neuron_5_mul_2_p <= Pix_68;
    10'd13:  neuron_5_mul_2_p <= Pix_69;
    10'd14:  neuron_5_mul_2_p <= Pix_70;
    10'd15:  neuron_5_mul_2_p <= Pix_71;
    10'd16:  neuron_5_mul_2_p <= Pix_72;
    10'd17:  neuron_5_mul_2_p <= Pix_73;
    10'd18:  neuron_5_mul_2_p <= Pix_74;
    10'd19:  neuron_5_mul_2_p <= Pix_75;
    10'd20:  neuron_5_mul_2_p <= Pix_76;
    10'd21:  neuron_5_mul_2_p <= Pix_77;
    10'd22:  neuron_5_mul_2_p <= Pix_78;
    10'd23:  neuron_5_mul_2_p <= Pix_79;
    10'd24:  neuron_5_mul_2_p <= Pix_80;
    10'd25:  neuron_5_mul_2_p <= Pix_81;
    10'd26:  neuron_5_mul_2_p <= Pix_82;
    10'd27:  neuron_5_mul_2_p <= Pix_83;
    default: neuron_5_mul_2_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_3_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_3_p <= Pix_84;
    10'd1:  neuron_5_mul_3_p <= Pix_85;
    10'd2:  neuron_5_mul_3_p <= Pix_86;
    10'd3:  neuron_5_mul_3_p <= Pix_87;
    10'd4:  neuron_5_mul_3_p <= Pix_88;
    10'd5:  neuron_5_mul_3_p <= Pix_89;
    10'd6:  neuron_5_mul_3_p <= Pix_90;
    10'd7:  neuron_5_mul_3_p <= Pix_91;
    10'd8:  neuron_5_mul_3_p <= Pix_92;
    10'd9:  neuron_5_mul_3_p <= Pix_93;
    10'd10:  neuron_5_mul_3_p <= Pix_94;
    10'd11:  neuron_5_mul_3_p <= Pix_95;
    10'd12:  neuron_5_mul_3_p <= Pix_96;
    10'd13:  neuron_5_mul_3_p <= Pix_97;
    10'd14:  neuron_5_mul_3_p <= Pix_98;
    10'd15:  neuron_5_mul_3_p <= Pix_99;
    10'd16:  neuron_5_mul_3_p <= Pix_100;
    10'd17:  neuron_5_mul_3_p <= Pix_101;
    10'd18:  neuron_5_mul_3_p <= Pix_102;
    10'd19:  neuron_5_mul_3_p <= Pix_103;
    10'd20:  neuron_5_mul_3_p <= Pix_104;
    10'd21:  neuron_5_mul_3_p <= Pix_105;
    10'd22:  neuron_5_mul_3_p <= Pix_106;
    10'd23:  neuron_5_mul_3_p <= Pix_107;
    10'd24:  neuron_5_mul_3_p <= Pix_108;
    10'd25:  neuron_5_mul_3_p <= Pix_109;
    10'd26:  neuron_5_mul_3_p <= Pix_110;
    10'd27:  neuron_5_mul_3_p <= Pix_111;
    default: neuron_5_mul_3_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_4_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_4_p <= Pix_112;
    10'd1:  neuron_5_mul_4_p <= Pix_113;
    10'd2:  neuron_5_mul_4_p <= Pix_114;
    10'd3:  neuron_5_mul_4_p <= Pix_115;
    10'd4:  neuron_5_mul_4_p <= Pix_116;
    10'd5:  neuron_5_mul_4_p <= Pix_117;
    10'd6:  neuron_5_mul_4_p <= Pix_118;
    10'd7:  neuron_5_mul_4_p <= Pix_119;
    10'd8:  neuron_5_mul_4_p <= Pix_120;
    10'd9:  neuron_5_mul_4_p <= Pix_121;
    10'd10:  neuron_5_mul_4_p <= Pix_122;
    10'd11:  neuron_5_mul_4_p <= Pix_123;
    10'd12:  neuron_5_mul_4_p <= Pix_124;
    10'd13:  neuron_5_mul_4_p <= Pix_125;
    10'd14:  neuron_5_mul_4_p <= Pix_126;
    10'd15:  neuron_5_mul_4_p <= Pix_127;
    10'd16:  neuron_5_mul_4_p <= Pix_128;
    10'd17:  neuron_5_mul_4_p <= Pix_129;
    10'd18:  neuron_5_mul_4_p <= Pix_130;
    10'd19:  neuron_5_mul_4_p <= Pix_131;
    10'd20:  neuron_5_mul_4_p <= Pix_132;
    10'd21:  neuron_5_mul_4_p <= Pix_133;
    10'd22:  neuron_5_mul_4_p <= Pix_134;
    10'd23:  neuron_5_mul_4_p <= Pix_135;
    10'd24:  neuron_5_mul_4_p <= Pix_136;
    10'd25:  neuron_5_mul_4_p <= Pix_137;
    10'd26:  neuron_5_mul_4_p <= Pix_138;
    10'd27:  neuron_5_mul_4_p <= Pix_139;
    default: neuron_5_mul_4_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_5_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_5_p <= Pix_140;
    10'd1:  neuron_5_mul_5_p <= Pix_141;
    10'd2:  neuron_5_mul_5_p <= Pix_142;
    10'd3:  neuron_5_mul_5_p <= Pix_143;
    10'd4:  neuron_5_mul_5_p <= Pix_144;
    10'd5:  neuron_5_mul_5_p <= Pix_145;
    10'd6:  neuron_5_mul_5_p <= Pix_146;
    10'd7:  neuron_5_mul_5_p <= Pix_147;
    10'd8:  neuron_5_mul_5_p <= Pix_148;
    10'd9:  neuron_5_mul_5_p <= Pix_149;
    10'd10:  neuron_5_mul_5_p <= Pix_150;
    10'd11:  neuron_5_mul_5_p <= Pix_151;
    10'd12:  neuron_5_mul_5_p <= Pix_152;
    10'd13:  neuron_5_mul_5_p <= Pix_153;
    10'd14:  neuron_5_mul_5_p <= Pix_154;
    10'd15:  neuron_5_mul_5_p <= Pix_155;
    10'd16:  neuron_5_mul_5_p <= Pix_156;
    10'd17:  neuron_5_mul_5_p <= Pix_157;
    10'd18:  neuron_5_mul_5_p <= Pix_158;
    10'd19:  neuron_5_mul_5_p <= Pix_159;
    10'd20:  neuron_5_mul_5_p <= Pix_160;
    10'd21:  neuron_5_mul_5_p <= Pix_161;
    10'd22:  neuron_5_mul_5_p <= Pix_162;
    10'd23:  neuron_5_mul_5_p <= Pix_163;
    10'd24:  neuron_5_mul_5_p <= Pix_164;
    10'd25:  neuron_5_mul_5_p <= Pix_165;
    10'd26:  neuron_5_mul_5_p <= Pix_166;
    10'd27:  neuron_5_mul_5_p <= Pix_167;
    default: neuron_5_mul_5_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_6_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_6_p <= Pix_168;
    10'd1:  neuron_5_mul_6_p <= Pix_169;
    10'd2:  neuron_5_mul_6_p <= Pix_170;
    10'd3:  neuron_5_mul_6_p <= Pix_171;
    10'd4:  neuron_5_mul_6_p <= Pix_172;
    10'd5:  neuron_5_mul_6_p <= Pix_173;
    10'd6:  neuron_5_mul_6_p <= Pix_174;
    10'd7:  neuron_5_mul_6_p <= Pix_175;
    10'd8:  neuron_5_mul_6_p <= Pix_176;
    10'd9:  neuron_5_mul_6_p <= Pix_177;
    10'd10:  neuron_5_mul_6_p <= Pix_178;
    10'd11:  neuron_5_mul_6_p <= Pix_179;
    10'd12:  neuron_5_mul_6_p <= Pix_180;
    10'd13:  neuron_5_mul_6_p <= Pix_181;
    10'd14:  neuron_5_mul_6_p <= Pix_182;
    10'd15:  neuron_5_mul_6_p <= Pix_183;
    10'd16:  neuron_5_mul_6_p <= Pix_184;
    10'd17:  neuron_5_mul_6_p <= Pix_185;
    10'd18:  neuron_5_mul_6_p <= Pix_186;
    10'd19:  neuron_5_mul_6_p <= Pix_187;
    10'd20:  neuron_5_mul_6_p <= Pix_188;
    10'd21:  neuron_5_mul_6_p <= Pix_189;
    10'd22:  neuron_5_mul_6_p <= Pix_190;
    10'd23:  neuron_5_mul_6_p <= Pix_191;
    10'd24:  neuron_5_mul_6_p <= Pix_192;
    10'd25:  neuron_5_mul_6_p <= Pix_193;
    10'd26:  neuron_5_mul_6_p <= Pix_194;
    10'd27:  neuron_5_mul_6_p <= Pix_195;
    default: neuron_5_mul_6_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_7_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_7_p <= Pix_196;
    10'd1:  neuron_5_mul_7_p <= Pix_197;
    10'd2:  neuron_5_mul_7_p <= Pix_198;
    10'd3:  neuron_5_mul_7_p <= Pix_199;
    10'd4:  neuron_5_mul_7_p <= Pix_200;
    10'd5:  neuron_5_mul_7_p <= Pix_201;
    10'd6:  neuron_5_mul_7_p <= Pix_202;
    10'd7:  neuron_5_mul_7_p <= Pix_203;
    10'd8:  neuron_5_mul_7_p <= Pix_204;
    10'd9:  neuron_5_mul_7_p <= Pix_205;
    10'd10:  neuron_5_mul_7_p <= Pix_206;
    10'd11:  neuron_5_mul_7_p <= Pix_207;
    10'd12:  neuron_5_mul_7_p <= Pix_208;
    10'd13:  neuron_5_mul_7_p <= Pix_209;
    10'd14:  neuron_5_mul_7_p <= Pix_210;
    10'd15:  neuron_5_mul_7_p <= Pix_211;
    10'd16:  neuron_5_mul_7_p <= Pix_212;
    10'd17:  neuron_5_mul_7_p <= Pix_213;
    10'd18:  neuron_5_mul_7_p <= Pix_214;
    10'd19:  neuron_5_mul_7_p <= Pix_215;
    10'd20:  neuron_5_mul_7_p <= Pix_216;
    10'd21:  neuron_5_mul_7_p <= Pix_217;
    10'd22:  neuron_5_mul_7_p <= Pix_218;
    10'd23:  neuron_5_mul_7_p <= Pix_219;
    10'd24:  neuron_5_mul_7_p <= Pix_220;
    10'd25:  neuron_5_mul_7_p <= Pix_221;
    10'd26:  neuron_5_mul_7_p <= Pix_222;
    10'd27:  neuron_5_mul_7_p <= Pix_223;
    default: neuron_5_mul_7_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_8_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_8_p <= Pix_224;
    10'd1:  neuron_5_mul_8_p <= Pix_225;
    10'd2:  neuron_5_mul_8_p <= Pix_226;
    10'd3:  neuron_5_mul_8_p <= Pix_227;
    10'd4:  neuron_5_mul_8_p <= Pix_228;
    10'd5:  neuron_5_mul_8_p <= Pix_229;
    10'd6:  neuron_5_mul_8_p <= Pix_230;
    10'd7:  neuron_5_mul_8_p <= Pix_231;
    10'd8:  neuron_5_mul_8_p <= Pix_232;
    10'd9:  neuron_5_mul_8_p <= Pix_233;
    10'd10:  neuron_5_mul_8_p <= Pix_234;
    10'd11:  neuron_5_mul_8_p <= Pix_235;
    10'd12:  neuron_5_mul_8_p <= Pix_236;
    10'd13:  neuron_5_mul_8_p <= Pix_237;
    10'd14:  neuron_5_mul_8_p <= Pix_238;
    10'd15:  neuron_5_mul_8_p <= Pix_239;
    10'd16:  neuron_5_mul_8_p <= Pix_240;
    10'd17:  neuron_5_mul_8_p <= Pix_241;
    10'd18:  neuron_5_mul_8_p <= Pix_242;
    10'd19:  neuron_5_mul_8_p <= Pix_243;
    10'd20:  neuron_5_mul_8_p <= Pix_244;
    10'd21:  neuron_5_mul_8_p <= Pix_245;
    10'd22:  neuron_5_mul_8_p <= Pix_246;
    10'd23:  neuron_5_mul_8_p <= Pix_247;
    10'd24:  neuron_5_mul_8_p <= Pix_248;
    10'd25:  neuron_5_mul_8_p <= Pix_249;
    10'd26:  neuron_5_mul_8_p <= Pix_250;
    10'd27:  neuron_5_mul_8_p <= Pix_251;
    default: neuron_5_mul_8_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_9_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_9_p <= Pix_252;
    10'd1:  neuron_5_mul_9_p <= Pix_253;
    10'd2:  neuron_5_mul_9_p <= Pix_254;
    10'd3:  neuron_5_mul_9_p <= Pix_255;
    10'd4:  neuron_5_mul_9_p <= Pix_256;
    10'd5:  neuron_5_mul_9_p <= Pix_257;
    10'd6:  neuron_5_mul_9_p <= Pix_258;
    10'd7:  neuron_5_mul_9_p <= Pix_259;
    10'd8:  neuron_5_mul_9_p <= Pix_260;
    10'd9:  neuron_5_mul_9_p <= Pix_261;
    10'd10:  neuron_5_mul_9_p <= Pix_262;
    10'd11:  neuron_5_mul_9_p <= Pix_263;
    10'd12:  neuron_5_mul_9_p <= Pix_264;
    10'd13:  neuron_5_mul_9_p <= Pix_265;
    10'd14:  neuron_5_mul_9_p <= Pix_266;
    10'd15:  neuron_5_mul_9_p <= Pix_267;
    10'd16:  neuron_5_mul_9_p <= Pix_268;
    10'd17:  neuron_5_mul_9_p <= Pix_269;
    10'd18:  neuron_5_mul_9_p <= Pix_270;
    10'd19:  neuron_5_mul_9_p <= Pix_271;
    10'd20:  neuron_5_mul_9_p <= Pix_272;
    10'd21:  neuron_5_mul_9_p <= Pix_273;
    10'd22:  neuron_5_mul_9_p <= Pix_274;
    10'd23:  neuron_5_mul_9_p <= Pix_275;
    10'd24:  neuron_5_mul_9_p <= Pix_276;
    10'd25:  neuron_5_mul_9_p <= Pix_277;
    10'd26:  neuron_5_mul_9_p <= Pix_278;
    10'd27:  neuron_5_mul_9_p <= Pix_279;
    default: neuron_5_mul_9_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_10_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_10_p <= Pix_280;
    10'd1:  neuron_5_mul_10_p <= Pix_281;
    10'd2:  neuron_5_mul_10_p <= Pix_282;
    10'd3:  neuron_5_mul_10_p <= Pix_283;
    10'd4:  neuron_5_mul_10_p <= Pix_284;
    10'd5:  neuron_5_mul_10_p <= Pix_285;
    10'd6:  neuron_5_mul_10_p <= Pix_286;
    10'd7:  neuron_5_mul_10_p <= Pix_287;
    10'd8:  neuron_5_mul_10_p <= Pix_288;
    10'd9:  neuron_5_mul_10_p <= Pix_289;
    10'd10:  neuron_5_mul_10_p <= Pix_290;
    10'd11:  neuron_5_mul_10_p <= Pix_291;
    10'd12:  neuron_5_mul_10_p <= Pix_292;
    10'd13:  neuron_5_mul_10_p <= Pix_293;
    10'd14:  neuron_5_mul_10_p <= Pix_294;
    10'd15:  neuron_5_mul_10_p <= Pix_295;
    10'd16:  neuron_5_mul_10_p <= Pix_296;
    10'd17:  neuron_5_mul_10_p <= Pix_297;
    10'd18:  neuron_5_mul_10_p <= Pix_298;
    10'd19:  neuron_5_mul_10_p <= Pix_299;
    10'd20:  neuron_5_mul_10_p <= Pix_300;
    10'd21:  neuron_5_mul_10_p <= Pix_301;
    10'd22:  neuron_5_mul_10_p <= Pix_302;
    10'd23:  neuron_5_mul_10_p <= Pix_303;
    10'd24:  neuron_5_mul_10_p <= Pix_304;
    10'd25:  neuron_5_mul_10_p <= Pix_305;
    10'd26:  neuron_5_mul_10_p <= Pix_306;
    10'd27:  neuron_5_mul_10_p <= Pix_307;
    default: neuron_5_mul_10_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_11_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_11_p <= Pix_308;
    10'd1:  neuron_5_mul_11_p <= Pix_309;
    10'd2:  neuron_5_mul_11_p <= Pix_310;
    10'd3:  neuron_5_mul_11_p <= Pix_311;
    10'd4:  neuron_5_mul_11_p <= Pix_312;
    10'd5:  neuron_5_mul_11_p <= Pix_313;
    10'd6:  neuron_5_mul_11_p <= Pix_314;
    10'd7:  neuron_5_mul_11_p <= Pix_315;
    10'd8:  neuron_5_mul_11_p <= Pix_316;
    10'd9:  neuron_5_mul_11_p <= Pix_317;
    10'd10:  neuron_5_mul_11_p <= Pix_318;
    10'd11:  neuron_5_mul_11_p <= Pix_319;
    10'd12:  neuron_5_mul_11_p <= Pix_320;
    10'd13:  neuron_5_mul_11_p <= Pix_321;
    10'd14:  neuron_5_mul_11_p <= Pix_322;
    10'd15:  neuron_5_mul_11_p <= Pix_323;
    10'd16:  neuron_5_mul_11_p <= Pix_324;
    10'd17:  neuron_5_mul_11_p <= Pix_325;
    10'd18:  neuron_5_mul_11_p <= Pix_326;
    10'd19:  neuron_5_mul_11_p <= Pix_327;
    10'd20:  neuron_5_mul_11_p <= Pix_328;
    10'd21:  neuron_5_mul_11_p <= Pix_329;
    10'd22:  neuron_5_mul_11_p <= Pix_330;
    10'd23:  neuron_5_mul_11_p <= Pix_331;
    10'd24:  neuron_5_mul_11_p <= Pix_332;
    10'd25:  neuron_5_mul_11_p <= Pix_333;
    10'd26:  neuron_5_mul_11_p <= Pix_334;
    10'd27:  neuron_5_mul_11_p <= Pix_335;
    default: neuron_5_mul_11_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_12_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_12_p <= Pix_336;
    10'd1:  neuron_5_mul_12_p <= Pix_337;
    10'd2:  neuron_5_mul_12_p <= Pix_338;
    10'd3:  neuron_5_mul_12_p <= Pix_339;
    10'd4:  neuron_5_mul_12_p <= Pix_340;
    10'd5:  neuron_5_mul_12_p <= Pix_341;
    10'd6:  neuron_5_mul_12_p <= Pix_342;
    10'd7:  neuron_5_mul_12_p <= Pix_343;
    10'd8:  neuron_5_mul_12_p <= Pix_344;
    10'd9:  neuron_5_mul_12_p <= Pix_345;
    10'd10:  neuron_5_mul_12_p <= Pix_346;
    10'd11:  neuron_5_mul_12_p <= Pix_347;
    10'd12:  neuron_5_mul_12_p <= Pix_348;
    10'd13:  neuron_5_mul_12_p <= Pix_349;
    10'd14:  neuron_5_mul_12_p <= Pix_350;
    10'd15:  neuron_5_mul_12_p <= Pix_351;
    10'd16:  neuron_5_mul_12_p <= Pix_352;
    10'd17:  neuron_5_mul_12_p <= Pix_353;
    10'd18:  neuron_5_mul_12_p <= Pix_354;
    10'd19:  neuron_5_mul_12_p <= Pix_355;
    10'd20:  neuron_5_mul_12_p <= Pix_356;
    10'd21:  neuron_5_mul_12_p <= Pix_357;
    10'd22:  neuron_5_mul_12_p <= Pix_358;
    10'd23:  neuron_5_mul_12_p <= Pix_359;
    10'd24:  neuron_5_mul_12_p <= Pix_360;
    10'd25:  neuron_5_mul_12_p <= Pix_361;
    10'd26:  neuron_5_mul_12_p <= Pix_362;
    10'd27:  neuron_5_mul_12_p <= Pix_363;
    default: neuron_5_mul_12_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_13_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_13_p <= Pix_364;
    10'd1:  neuron_5_mul_13_p <= Pix_365;
    10'd2:  neuron_5_mul_13_p <= Pix_366;
    10'd3:  neuron_5_mul_13_p <= Pix_367;
    10'd4:  neuron_5_mul_13_p <= Pix_368;
    10'd5:  neuron_5_mul_13_p <= Pix_369;
    10'd6:  neuron_5_mul_13_p <= Pix_370;
    10'd7:  neuron_5_mul_13_p <= Pix_371;
    10'd8:  neuron_5_mul_13_p <= Pix_372;
    10'd9:  neuron_5_mul_13_p <= Pix_373;
    10'd10:  neuron_5_mul_13_p <= Pix_374;
    10'd11:  neuron_5_mul_13_p <= Pix_375;
    10'd12:  neuron_5_mul_13_p <= Pix_376;
    10'd13:  neuron_5_mul_13_p <= Pix_377;
    10'd14:  neuron_5_mul_13_p <= Pix_378;
    10'd15:  neuron_5_mul_13_p <= Pix_379;
    10'd16:  neuron_5_mul_13_p <= Pix_380;
    10'd17:  neuron_5_mul_13_p <= Pix_381;
    10'd18:  neuron_5_mul_13_p <= Pix_382;
    10'd19:  neuron_5_mul_13_p <= Pix_383;
    10'd20:  neuron_5_mul_13_p <= Pix_384;
    10'd21:  neuron_5_mul_13_p <= Pix_385;
    10'd22:  neuron_5_mul_13_p <= Pix_386;
    10'd23:  neuron_5_mul_13_p <= Pix_387;
    10'd24:  neuron_5_mul_13_p <= Pix_388;
    10'd25:  neuron_5_mul_13_p <= Pix_389;
    10'd26:  neuron_5_mul_13_p <= Pix_390;
    10'd27:  neuron_5_mul_13_p <= Pix_391;
    default: neuron_5_mul_13_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_14_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_14_p <= Pix_392;
    10'd1:  neuron_5_mul_14_p <= Pix_393;
    10'd2:  neuron_5_mul_14_p <= Pix_394;
    10'd3:  neuron_5_mul_14_p <= Pix_395;
    10'd4:  neuron_5_mul_14_p <= Pix_396;
    10'd5:  neuron_5_mul_14_p <= Pix_397;
    10'd6:  neuron_5_mul_14_p <= Pix_398;
    10'd7:  neuron_5_mul_14_p <= Pix_399;
    10'd8:  neuron_5_mul_14_p <= Pix_400;
    10'd9:  neuron_5_mul_14_p <= Pix_401;
    10'd10:  neuron_5_mul_14_p <= Pix_402;
    10'd11:  neuron_5_mul_14_p <= Pix_403;
    10'd12:  neuron_5_mul_14_p <= Pix_404;
    10'd13:  neuron_5_mul_14_p <= Pix_405;
    10'd14:  neuron_5_mul_14_p <= Pix_406;
    10'd15:  neuron_5_mul_14_p <= Pix_407;
    10'd16:  neuron_5_mul_14_p <= Pix_408;
    10'd17:  neuron_5_mul_14_p <= Pix_409;
    10'd18:  neuron_5_mul_14_p <= Pix_410;
    10'd19:  neuron_5_mul_14_p <= Pix_411;
    10'd20:  neuron_5_mul_14_p <= Pix_412;
    10'd21:  neuron_5_mul_14_p <= Pix_413;
    10'd22:  neuron_5_mul_14_p <= Pix_414;
    10'd23:  neuron_5_mul_14_p <= Pix_415;
    10'd24:  neuron_5_mul_14_p <= Pix_416;
    10'd25:  neuron_5_mul_14_p <= Pix_417;
    10'd26:  neuron_5_mul_14_p <= Pix_418;
    10'd27:  neuron_5_mul_14_p <= Pix_419;
    default: neuron_5_mul_14_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_15_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_15_p <= Pix_420;
    10'd1:  neuron_5_mul_15_p <= Pix_421;
    10'd2:  neuron_5_mul_15_p <= Pix_422;
    10'd3:  neuron_5_mul_15_p <= Pix_423;
    10'd4:  neuron_5_mul_15_p <= Pix_424;
    10'd5:  neuron_5_mul_15_p <= Pix_425;
    10'd6:  neuron_5_mul_15_p <= Pix_426;
    10'd7:  neuron_5_mul_15_p <= Pix_427;
    10'd8:  neuron_5_mul_15_p <= Pix_428;
    10'd9:  neuron_5_mul_15_p <= Pix_429;
    10'd10:  neuron_5_mul_15_p <= Pix_430;
    10'd11:  neuron_5_mul_15_p <= Pix_431;
    10'd12:  neuron_5_mul_15_p <= Pix_432;
    10'd13:  neuron_5_mul_15_p <= Pix_433;
    10'd14:  neuron_5_mul_15_p <= Pix_434;
    10'd15:  neuron_5_mul_15_p <= Pix_435;
    10'd16:  neuron_5_mul_15_p <= Pix_436;
    10'd17:  neuron_5_mul_15_p <= Pix_437;
    10'd18:  neuron_5_mul_15_p <= Pix_438;
    10'd19:  neuron_5_mul_15_p <= Pix_439;
    10'd20:  neuron_5_mul_15_p <= Pix_440;
    10'd21:  neuron_5_mul_15_p <= Pix_441;
    10'd22:  neuron_5_mul_15_p <= Pix_442;
    10'd23:  neuron_5_mul_15_p <= Pix_443;
    10'd24:  neuron_5_mul_15_p <= Pix_444;
    10'd25:  neuron_5_mul_15_p <= Pix_445;
    10'd26:  neuron_5_mul_15_p <= Pix_446;
    10'd27:  neuron_5_mul_15_p <= Pix_447;
    default: neuron_5_mul_15_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_16_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_16_p <= Pix_448;
    10'd1:  neuron_5_mul_16_p <= Pix_449;
    10'd2:  neuron_5_mul_16_p <= Pix_450;
    10'd3:  neuron_5_mul_16_p <= Pix_451;
    10'd4:  neuron_5_mul_16_p <= Pix_452;
    10'd5:  neuron_5_mul_16_p <= Pix_453;
    10'd6:  neuron_5_mul_16_p <= Pix_454;
    10'd7:  neuron_5_mul_16_p <= Pix_455;
    10'd8:  neuron_5_mul_16_p <= Pix_456;
    10'd9:  neuron_5_mul_16_p <= Pix_457;
    10'd10:  neuron_5_mul_16_p <= Pix_458;
    10'd11:  neuron_5_mul_16_p <= Pix_459;
    10'd12:  neuron_5_mul_16_p <= Pix_460;
    10'd13:  neuron_5_mul_16_p <= Pix_461;
    10'd14:  neuron_5_mul_16_p <= Pix_462;
    10'd15:  neuron_5_mul_16_p <= Pix_463;
    10'd16:  neuron_5_mul_16_p <= Pix_464;
    10'd17:  neuron_5_mul_16_p <= Pix_465;
    10'd18:  neuron_5_mul_16_p <= Pix_466;
    10'd19:  neuron_5_mul_16_p <= Pix_467;
    10'd20:  neuron_5_mul_16_p <= Pix_468;
    10'd21:  neuron_5_mul_16_p <= Pix_469;
    10'd22:  neuron_5_mul_16_p <= Pix_470;
    10'd23:  neuron_5_mul_16_p <= Pix_471;
    10'd24:  neuron_5_mul_16_p <= Pix_472;
    10'd25:  neuron_5_mul_16_p <= Pix_473;
    10'd26:  neuron_5_mul_16_p <= Pix_474;
    10'd27:  neuron_5_mul_16_p <= Pix_475;
    default: neuron_5_mul_16_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_17_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_17_p <= Pix_476;
    10'd1:  neuron_5_mul_17_p <= Pix_477;
    10'd2:  neuron_5_mul_17_p <= Pix_478;
    10'd3:  neuron_5_mul_17_p <= Pix_479;
    10'd4:  neuron_5_mul_17_p <= Pix_480;
    10'd5:  neuron_5_mul_17_p <= Pix_481;
    10'd6:  neuron_5_mul_17_p <= Pix_482;
    10'd7:  neuron_5_mul_17_p <= Pix_483;
    10'd8:  neuron_5_mul_17_p <= Pix_484;
    10'd9:  neuron_5_mul_17_p <= Pix_485;
    10'd10:  neuron_5_mul_17_p <= Pix_486;
    10'd11:  neuron_5_mul_17_p <= Pix_487;
    10'd12:  neuron_5_mul_17_p <= Pix_488;
    10'd13:  neuron_5_mul_17_p <= Pix_489;
    10'd14:  neuron_5_mul_17_p <= Pix_490;
    10'd15:  neuron_5_mul_17_p <= Pix_491;
    10'd16:  neuron_5_mul_17_p <= Pix_492;
    10'd17:  neuron_5_mul_17_p <= Pix_493;
    10'd18:  neuron_5_mul_17_p <= Pix_494;
    10'd19:  neuron_5_mul_17_p <= Pix_495;
    10'd20:  neuron_5_mul_17_p <= Pix_496;
    10'd21:  neuron_5_mul_17_p <= Pix_497;
    10'd22:  neuron_5_mul_17_p <= Pix_498;
    10'd23:  neuron_5_mul_17_p <= Pix_499;
    10'd24:  neuron_5_mul_17_p <= Pix_500;
    10'd25:  neuron_5_mul_17_p <= Pix_501;
    10'd26:  neuron_5_mul_17_p <= Pix_502;
    10'd27:  neuron_5_mul_17_p <= Pix_503;
    default: neuron_5_mul_17_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_18_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_18_p <= Pix_504;
    10'd1:  neuron_5_mul_18_p <= Pix_505;
    10'd2:  neuron_5_mul_18_p <= Pix_506;
    10'd3:  neuron_5_mul_18_p <= Pix_507;
    10'd4:  neuron_5_mul_18_p <= Pix_508;
    10'd5:  neuron_5_mul_18_p <= Pix_509;
    10'd6:  neuron_5_mul_18_p <= Pix_510;
    10'd7:  neuron_5_mul_18_p <= Pix_511;
    10'd8:  neuron_5_mul_18_p <= Pix_512;
    10'd9:  neuron_5_mul_18_p <= Pix_513;
    10'd10:  neuron_5_mul_18_p <= Pix_514;
    10'd11:  neuron_5_mul_18_p <= Pix_515;
    10'd12:  neuron_5_mul_18_p <= Pix_516;
    10'd13:  neuron_5_mul_18_p <= Pix_517;
    10'd14:  neuron_5_mul_18_p <= Pix_518;
    10'd15:  neuron_5_mul_18_p <= Pix_519;
    10'd16:  neuron_5_mul_18_p <= Pix_520;
    10'd17:  neuron_5_mul_18_p <= Pix_521;
    10'd18:  neuron_5_mul_18_p <= Pix_522;
    10'd19:  neuron_5_mul_18_p <= Pix_523;
    10'd20:  neuron_5_mul_18_p <= Pix_524;
    10'd21:  neuron_5_mul_18_p <= Pix_525;
    10'd22:  neuron_5_mul_18_p <= Pix_526;
    10'd23:  neuron_5_mul_18_p <= Pix_527;
    10'd24:  neuron_5_mul_18_p <= Pix_528;
    10'd25:  neuron_5_mul_18_p <= Pix_529;
    10'd26:  neuron_5_mul_18_p <= Pix_530;
    10'd27:  neuron_5_mul_18_p <= Pix_531;
    default: neuron_5_mul_18_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_19_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_19_p <= Pix_532;
    10'd1:  neuron_5_mul_19_p <= Pix_533;
    10'd2:  neuron_5_mul_19_p <= Pix_534;
    10'd3:  neuron_5_mul_19_p <= Pix_535;
    10'd4:  neuron_5_mul_19_p <= Pix_536;
    10'd5:  neuron_5_mul_19_p <= Pix_537;
    10'd6:  neuron_5_mul_19_p <= Pix_538;
    10'd7:  neuron_5_mul_19_p <= Pix_539;
    10'd8:  neuron_5_mul_19_p <= Pix_540;
    10'd9:  neuron_5_mul_19_p <= Pix_541;
    10'd10:  neuron_5_mul_19_p <= Pix_542;
    10'd11:  neuron_5_mul_19_p <= Pix_543;
    10'd12:  neuron_5_mul_19_p <= Pix_544;
    10'd13:  neuron_5_mul_19_p <= Pix_545;
    10'd14:  neuron_5_mul_19_p <= Pix_546;
    10'd15:  neuron_5_mul_19_p <= Pix_547;
    10'd16:  neuron_5_mul_19_p <= Pix_548;
    10'd17:  neuron_5_mul_19_p <= Pix_549;
    10'd18:  neuron_5_mul_19_p <= Pix_550;
    10'd19:  neuron_5_mul_19_p <= Pix_551;
    10'd20:  neuron_5_mul_19_p <= Pix_552;
    10'd21:  neuron_5_mul_19_p <= Pix_553;
    10'd22:  neuron_5_mul_19_p <= Pix_554;
    10'd23:  neuron_5_mul_19_p <= Pix_555;
    10'd24:  neuron_5_mul_19_p <= Pix_556;
    10'd25:  neuron_5_mul_19_p <= Pix_557;
    10'd26:  neuron_5_mul_19_p <= Pix_558;
    10'd27:  neuron_5_mul_19_p <= Pix_559;
    default: neuron_5_mul_19_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_20_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_20_p <= Pix_560;
    10'd1:  neuron_5_mul_20_p <= Pix_561;
    10'd2:  neuron_5_mul_20_p <= Pix_562;
    10'd3:  neuron_5_mul_20_p <= Pix_563;
    10'd4:  neuron_5_mul_20_p <= Pix_564;
    10'd5:  neuron_5_mul_20_p <= Pix_565;
    10'd6:  neuron_5_mul_20_p <= Pix_566;
    10'd7:  neuron_5_mul_20_p <= Pix_567;
    10'd8:  neuron_5_mul_20_p <= Pix_568;
    10'd9:  neuron_5_mul_20_p <= Pix_569;
    10'd10:  neuron_5_mul_20_p <= Pix_570;
    10'd11:  neuron_5_mul_20_p <= Pix_571;
    10'd12:  neuron_5_mul_20_p <= Pix_572;
    10'd13:  neuron_5_mul_20_p <= Pix_573;
    10'd14:  neuron_5_mul_20_p <= Pix_574;
    10'd15:  neuron_5_mul_20_p <= Pix_575;
    10'd16:  neuron_5_mul_20_p <= Pix_576;
    10'd17:  neuron_5_mul_20_p <= Pix_577;
    10'd18:  neuron_5_mul_20_p <= Pix_578;
    10'd19:  neuron_5_mul_20_p <= Pix_579;
    10'd20:  neuron_5_mul_20_p <= Pix_580;
    10'd21:  neuron_5_mul_20_p <= Pix_581;
    10'd22:  neuron_5_mul_20_p <= Pix_582;
    10'd23:  neuron_5_mul_20_p <= Pix_583;
    10'd24:  neuron_5_mul_20_p <= Pix_584;
    10'd25:  neuron_5_mul_20_p <= Pix_585;
    10'd26:  neuron_5_mul_20_p <= Pix_586;
    10'd27:  neuron_5_mul_20_p <= Pix_587;
    default: neuron_5_mul_20_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_21_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_21_p <= Pix_588;
    10'd1:  neuron_5_mul_21_p <= Pix_589;
    10'd2:  neuron_5_mul_21_p <= Pix_590;
    10'd3:  neuron_5_mul_21_p <= Pix_591;
    10'd4:  neuron_5_mul_21_p <= Pix_592;
    10'd5:  neuron_5_mul_21_p <= Pix_593;
    10'd6:  neuron_5_mul_21_p <= Pix_594;
    10'd7:  neuron_5_mul_21_p <= Pix_595;
    10'd8:  neuron_5_mul_21_p <= Pix_596;
    10'd9:  neuron_5_mul_21_p <= Pix_597;
    10'd10:  neuron_5_mul_21_p <= Pix_598;
    10'd11:  neuron_5_mul_21_p <= Pix_599;
    10'd12:  neuron_5_mul_21_p <= Pix_600;
    10'd13:  neuron_5_mul_21_p <= Pix_601;
    10'd14:  neuron_5_mul_21_p <= Pix_602;
    10'd15:  neuron_5_mul_21_p <= Pix_603;
    10'd16:  neuron_5_mul_21_p <= Pix_604;
    10'd17:  neuron_5_mul_21_p <= Pix_605;
    10'd18:  neuron_5_mul_21_p <= Pix_606;
    10'd19:  neuron_5_mul_21_p <= Pix_607;
    10'd20:  neuron_5_mul_21_p <= Pix_608;
    10'd21:  neuron_5_mul_21_p <= Pix_609;
    10'd22:  neuron_5_mul_21_p <= Pix_610;
    10'd23:  neuron_5_mul_21_p <= Pix_611;
    10'd24:  neuron_5_mul_21_p <= Pix_612;
    10'd25:  neuron_5_mul_21_p <= Pix_613;
    10'd26:  neuron_5_mul_21_p <= Pix_614;
    10'd27:  neuron_5_mul_21_p <= Pix_615;
    default: neuron_5_mul_21_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_22_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_22_p <= Pix_616;
    10'd1:  neuron_5_mul_22_p <= Pix_617;
    10'd2:  neuron_5_mul_22_p <= Pix_618;
    10'd3:  neuron_5_mul_22_p <= Pix_619;
    10'd4:  neuron_5_mul_22_p <= Pix_620;
    10'd5:  neuron_5_mul_22_p <= Pix_621;
    10'd6:  neuron_5_mul_22_p <= Pix_622;
    10'd7:  neuron_5_mul_22_p <= Pix_623;
    10'd8:  neuron_5_mul_22_p <= Pix_624;
    10'd9:  neuron_5_mul_22_p <= Pix_625;
    10'd10:  neuron_5_mul_22_p <= Pix_626;
    10'd11:  neuron_5_mul_22_p <= Pix_627;
    10'd12:  neuron_5_mul_22_p <= Pix_628;
    10'd13:  neuron_5_mul_22_p <= Pix_629;
    10'd14:  neuron_5_mul_22_p <= Pix_630;
    10'd15:  neuron_5_mul_22_p <= Pix_631;
    10'd16:  neuron_5_mul_22_p <= Pix_632;
    10'd17:  neuron_5_mul_22_p <= Pix_633;
    10'd18:  neuron_5_mul_22_p <= Pix_634;
    10'd19:  neuron_5_mul_22_p <= Pix_635;
    10'd20:  neuron_5_mul_22_p <= Pix_636;
    10'd21:  neuron_5_mul_22_p <= Pix_637;
    10'd22:  neuron_5_mul_22_p <= Pix_638;
    10'd23:  neuron_5_mul_22_p <= Pix_639;
    10'd24:  neuron_5_mul_22_p <= Pix_640;
    10'd25:  neuron_5_mul_22_p <= Pix_641;
    10'd26:  neuron_5_mul_22_p <= Pix_642;
    10'd27:  neuron_5_mul_22_p <= Pix_643;
    default: neuron_5_mul_22_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_23_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_23_p <= Pix_644;
    10'd1:  neuron_5_mul_23_p <= Pix_645;
    10'd2:  neuron_5_mul_23_p <= Pix_646;
    10'd3:  neuron_5_mul_23_p <= Pix_647;
    10'd4:  neuron_5_mul_23_p <= Pix_648;
    10'd5:  neuron_5_mul_23_p <= Pix_649;
    10'd6:  neuron_5_mul_23_p <= Pix_650;
    10'd7:  neuron_5_mul_23_p <= Pix_651;
    10'd8:  neuron_5_mul_23_p <= Pix_652;
    10'd9:  neuron_5_mul_23_p <= Pix_653;
    10'd10:  neuron_5_mul_23_p <= Pix_654;
    10'd11:  neuron_5_mul_23_p <= Pix_655;
    10'd12:  neuron_5_mul_23_p <= Pix_656;
    10'd13:  neuron_5_mul_23_p <= Pix_657;
    10'd14:  neuron_5_mul_23_p <= Pix_658;
    10'd15:  neuron_5_mul_23_p <= Pix_659;
    10'd16:  neuron_5_mul_23_p <= Pix_660;
    10'd17:  neuron_5_mul_23_p <= Pix_661;
    10'd18:  neuron_5_mul_23_p <= Pix_662;
    10'd19:  neuron_5_mul_23_p <= Pix_663;
    10'd20:  neuron_5_mul_23_p <= Pix_664;
    10'd21:  neuron_5_mul_23_p <= Pix_665;
    10'd22:  neuron_5_mul_23_p <= Pix_666;
    10'd23:  neuron_5_mul_23_p <= Pix_667;
    10'd24:  neuron_5_mul_23_p <= Pix_668;
    10'd25:  neuron_5_mul_23_p <= Pix_669;
    10'd26:  neuron_5_mul_23_p <= Pix_670;
    10'd27:  neuron_5_mul_23_p <= Pix_671;
    default: neuron_5_mul_23_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_24_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_24_p <= Pix_672;
    10'd1:  neuron_5_mul_24_p <= Pix_673;
    10'd2:  neuron_5_mul_24_p <= Pix_674;
    10'd3:  neuron_5_mul_24_p <= Pix_675;
    10'd4:  neuron_5_mul_24_p <= Pix_676;
    10'd5:  neuron_5_mul_24_p <= Pix_677;
    10'd6:  neuron_5_mul_24_p <= Pix_678;
    10'd7:  neuron_5_mul_24_p <= Pix_679;
    10'd8:  neuron_5_mul_24_p <= Pix_680;
    10'd9:  neuron_5_mul_24_p <= Pix_681;
    10'd10:  neuron_5_mul_24_p <= Pix_682;
    10'd11:  neuron_5_mul_24_p <= Pix_683;
    10'd12:  neuron_5_mul_24_p <= Pix_684;
    10'd13:  neuron_5_mul_24_p <= Pix_685;
    10'd14:  neuron_5_mul_24_p <= Pix_686;
    10'd15:  neuron_5_mul_24_p <= Pix_687;
    10'd16:  neuron_5_mul_24_p <= Pix_688;
    10'd17:  neuron_5_mul_24_p <= Pix_689;
    10'd18:  neuron_5_mul_24_p <= Pix_690;
    10'd19:  neuron_5_mul_24_p <= Pix_691;
    10'd20:  neuron_5_mul_24_p <= Pix_692;
    10'd21:  neuron_5_mul_24_p <= Pix_693;
    10'd22:  neuron_5_mul_24_p <= Pix_694;
    10'd23:  neuron_5_mul_24_p <= Pix_695;
    10'd24:  neuron_5_mul_24_p <= Pix_696;
    10'd25:  neuron_5_mul_24_p <= Pix_697;
    10'd26:  neuron_5_mul_24_p <= Pix_698;
    10'd27:  neuron_5_mul_24_p <= Pix_699;
    default: neuron_5_mul_24_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_25_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_25_p <= Pix_700;
    10'd1:  neuron_5_mul_25_p <= Pix_701;
    10'd2:  neuron_5_mul_25_p <= Pix_702;
    10'd3:  neuron_5_mul_25_p <= Pix_703;
    10'd4:  neuron_5_mul_25_p <= Pix_704;
    10'd5:  neuron_5_mul_25_p <= Pix_705;
    10'd6:  neuron_5_mul_25_p <= Pix_706;
    10'd7:  neuron_5_mul_25_p <= Pix_707;
    10'd8:  neuron_5_mul_25_p <= Pix_708;
    10'd9:  neuron_5_mul_25_p <= Pix_709;
    10'd10:  neuron_5_mul_25_p <= Pix_710;
    10'd11:  neuron_5_mul_25_p <= Pix_711;
    10'd12:  neuron_5_mul_25_p <= Pix_712;
    10'd13:  neuron_5_mul_25_p <= Pix_713;
    10'd14:  neuron_5_mul_25_p <= Pix_714;
    10'd15:  neuron_5_mul_25_p <= Pix_715;
    10'd16:  neuron_5_mul_25_p <= Pix_716;
    10'd17:  neuron_5_mul_25_p <= Pix_717;
    10'd18:  neuron_5_mul_25_p <= Pix_718;
    10'd19:  neuron_5_mul_25_p <= Pix_719;
    10'd20:  neuron_5_mul_25_p <= Pix_720;
    10'd21:  neuron_5_mul_25_p <= Pix_721;
    10'd22:  neuron_5_mul_25_p <= Pix_722;
    10'd23:  neuron_5_mul_25_p <= Pix_723;
    10'd24:  neuron_5_mul_25_p <= Pix_724;
    10'd25:  neuron_5_mul_25_p <= Pix_725;
    10'd26:  neuron_5_mul_25_p <= Pix_726;
    10'd27:  neuron_5_mul_25_p <= Pix_727;
    default: neuron_5_mul_25_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_26_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_26_p <= Pix_728;
    10'd1:  neuron_5_mul_26_p <= Pix_729;
    10'd2:  neuron_5_mul_26_p <= Pix_730;
    10'd3:  neuron_5_mul_26_p <= Pix_731;
    10'd4:  neuron_5_mul_26_p <= Pix_732;
    10'd5:  neuron_5_mul_26_p <= Pix_733;
    10'd6:  neuron_5_mul_26_p <= Pix_734;
    10'd7:  neuron_5_mul_26_p <= Pix_735;
    10'd8:  neuron_5_mul_26_p <= Pix_736;
    10'd9:  neuron_5_mul_26_p <= Pix_737;
    10'd10:  neuron_5_mul_26_p <= Pix_738;
    10'd11:  neuron_5_mul_26_p <= Pix_739;
    10'd12:  neuron_5_mul_26_p <= Pix_740;
    10'd13:  neuron_5_mul_26_p <= Pix_741;
    10'd14:  neuron_5_mul_26_p <= Pix_742;
    10'd15:  neuron_5_mul_26_p <= Pix_743;
    10'd16:  neuron_5_mul_26_p <= Pix_744;
    10'd17:  neuron_5_mul_26_p <= Pix_745;
    10'd18:  neuron_5_mul_26_p <= Pix_746;
    10'd19:  neuron_5_mul_26_p <= Pix_747;
    10'd20:  neuron_5_mul_26_p <= Pix_748;
    10'd21:  neuron_5_mul_26_p <= Pix_749;
    10'd22:  neuron_5_mul_26_p <= Pix_750;
    10'd23:  neuron_5_mul_26_p <= Pix_751;
    10'd24:  neuron_5_mul_26_p <= Pix_752;
    10'd25:  neuron_5_mul_26_p <= Pix_753;
    10'd26:  neuron_5_mul_26_p <= Pix_754;
    10'd27:  neuron_5_mul_26_p <= Pix_755;
    default: neuron_5_mul_26_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_5_mul_27_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_5_mul_27_p <= Pix_756;
    10'd1:  neuron_5_mul_27_p <= Pix_757;
    10'd2:  neuron_5_mul_27_p <= Pix_758;
    10'd3:  neuron_5_mul_27_p <= Pix_759;
    10'd4:  neuron_5_mul_27_p <= Pix_760;
    10'd5:  neuron_5_mul_27_p <= Pix_761;
    10'd6:  neuron_5_mul_27_p <= Pix_762;
    10'd7:  neuron_5_mul_27_p <= Pix_763;
    10'd8:  neuron_5_mul_27_p <= Pix_764;
    10'd9:  neuron_5_mul_27_p <= Pix_765;
    10'd10:  neuron_5_mul_27_p <= Pix_766;
    10'd11:  neuron_5_mul_27_p <= Pix_767;
    10'd12:  neuron_5_mul_27_p <= Pix_768;
    10'd13:  neuron_5_mul_27_p <= Pix_769;
    10'd14:  neuron_5_mul_27_p <= Pix_770;
    10'd15:  neuron_5_mul_27_p <= Pix_771;
    10'd16:  neuron_5_mul_27_p <= Pix_772;
    10'd17:  neuron_5_mul_27_p <= Pix_773;
    10'd18:  neuron_5_mul_27_p <= Pix_774;
    10'd19:  neuron_5_mul_27_p <= Pix_775;
    10'd20:  neuron_5_mul_27_p <= Pix_776;
    10'd21:  neuron_5_mul_27_p <= Pix_777;
    10'd22:  neuron_5_mul_27_p <= Pix_778;
    10'd23:  neuron_5_mul_27_p <= Pix_779;
    10'd24:  neuron_5_mul_27_p <= Pix_780;
    10'd25:  neuron_5_mul_27_p <= Pix_781;
    10'd26:  neuron_5_mul_27_p <= Pix_782;
    10'd27:  neuron_5_mul_27_p <= Pix_783;
    default: neuron_5_mul_27_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_0_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_0_p <= Pix_0;
    10'd1:  neuron_6_mul_0_p <= Pix_1;
    10'd2:  neuron_6_mul_0_p <= Pix_2;
    10'd3:  neuron_6_mul_0_p <= Pix_3;
    10'd4:  neuron_6_mul_0_p <= Pix_4;
    10'd5:  neuron_6_mul_0_p <= Pix_5;
    10'd6:  neuron_6_mul_0_p <= Pix_6;
    10'd7:  neuron_6_mul_0_p <= Pix_7;
    10'd8:  neuron_6_mul_0_p <= Pix_8;
    10'd9:  neuron_6_mul_0_p <= Pix_9;
    10'd10:  neuron_6_mul_0_p <= Pix_10;
    10'd11:  neuron_6_mul_0_p <= Pix_11;
    10'd12:  neuron_6_mul_0_p <= Pix_12;
    10'd13:  neuron_6_mul_0_p <= Pix_13;
    10'd14:  neuron_6_mul_0_p <= Pix_14;
    10'd15:  neuron_6_mul_0_p <= Pix_15;
    10'd16:  neuron_6_mul_0_p <= Pix_16;
    10'd17:  neuron_6_mul_0_p <= Pix_17;
    10'd18:  neuron_6_mul_0_p <= Pix_18;
    10'd19:  neuron_6_mul_0_p <= Pix_19;
    10'd20:  neuron_6_mul_0_p <= Pix_20;
    10'd21:  neuron_6_mul_0_p <= Pix_21;
    10'd22:  neuron_6_mul_0_p <= Pix_22;
    10'd23:  neuron_6_mul_0_p <= Pix_23;
    10'd24:  neuron_6_mul_0_p <= Pix_24;
    10'd25:  neuron_6_mul_0_p <= Pix_25;
    10'd26:  neuron_6_mul_0_p <= Pix_26;
    10'd27:  neuron_6_mul_0_p <= Pix_27;
    default: neuron_6_mul_0_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_1_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_1_p <= Pix_28;
    10'd1:  neuron_6_mul_1_p <= Pix_29;
    10'd2:  neuron_6_mul_1_p <= Pix_30;
    10'd3:  neuron_6_mul_1_p <= Pix_31;
    10'd4:  neuron_6_mul_1_p <= Pix_32;
    10'd5:  neuron_6_mul_1_p <= Pix_33;
    10'd6:  neuron_6_mul_1_p <= Pix_34;
    10'd7:  neuron_6_mul_1_p <= Pix_35;
    10'd8:  neuron_6_mul_1_p <= Pix_36;
    10'd9:  neuron_6_mul_1_p <= Pix_37;
    10'd10:  neuron_6_mul_1_p <= Pix_38;
    10'd11:  neuron_6_mul_1_p <= Pix_39;
    10'd12:  neuron_6_mul_1_p <= Pix_40;
    10'd13:  neuron_6_mul_1_p <= Pix_41;
    10'd14:  neuron_6_mul_1_p <= Pix_42;
    10'd15:  neuron_6_mul_1_p <= Pix_43;
    10'd16:  neuron_6_mul_1_p <= Pix_44;
    10'd17:  neuron_6_mul_1_p <= Pix_45;
    10'd18:  neuron_6_mul_1_p <= Pix_46;
    10'd19:  neuron_6_mul_1_p <= Pix_47;
    10'd20:  neuron_6_mul_1_p <= Pix_48;
    10'd21:  neuron_6_mul_1_p <= Pix_49;
    10'd22:  neuron_6_mul_1_p <= Pix_50;
    10'd23:  neuron_6_mul_1_p <= Pix_51;
    10'd24:  neuron_6_mul_1_p <= Pix_52;
    10'd25:  neuron_6_mul_1_p <= Pix_53;
    10'd26:  neuron_6_mul_1_p <= Pix_54;
    10'd27:  neuron_6_mul_1_p <= Pix_55;
    default: neuron_6_mul_1_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_2_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_2_p <= Pix_56;
    10'd1:  neuron_6_mul_2_p <= Pix_57;
    10'd2:  neuron_6_mul_2_p <= Pix_58;
    10'd3:  neuron_6_mul_2_p <= Pix_59;
    10'd4:  neuron_6_mul_2_p <= Pix_60;
    10'd5:  neuron_6_mul_2_p <= Pix_61;
    10'd6:  neuron_6_mul_2_p <= Pix_62;
    10'd7:  neuron_6_mul_2_p <= Pix_63;
    10'd8:  neuron_6_mul_2_p <= Pix_64;
    10'd9:  neuron_6_mul_2_p <= Pix_65;
    10'd10:  neuron_6_mul_2_p <= Pix_66;
    10'd11:  neuron_6_mul_2_p <= Pix_67;
    10'd12:  neuron_6_mul_2_p <= Pix_68;
    10'd13:  neuron_6_mul_2_p <= Pix_69;
    10'd14:  neuron_6_mul_2_p <= Pix_70;
    10'd15:  neuron_6_mul_2_p <= Pix_71;
    10'd16:  neuron_6_mul_2_p <= Pix_72;
    10'd17:  neuron_6_mul_2_p <= Pix_73;
    10'd18:  neuron_6_mul_2_p <= Pix_74;
    10'd19:  neuron_6_mul_2_p <= Pix_75;
    10'd20:  neuron_6_mul_2_p <= Pix_76;
    10'd21:  neuron_6_mul_2_p <= Pix_77;
    10'd22:  neuron_6_mul_2_p <= Pix_78;
    10'd23:  neuron_6_mul_2_p <= Pix_79;
    10'd24:  neuron_6_mul_2_p <= Pix_80;
    10'd25:  neuron_6_mul_2_p <= Pix_81;
    10'd26:  neuron_6_mul_2_p <= Pix_82;
    10'd27:  neuron_6_mul_2_p <= Pix_83;
    default: neuron_6_mul_2_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_3_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_3_p <= Pix_84;
    10'd1:  neuron_6_mul_3_p <= Pix_85;
    10'd2:  neuron_6_mul_3_p <= Pix_86;
    10'd3:  neuron_6_mul_3_p <= Pix_87;
    10'd4:  neuron_6_mul_3_p <= Pix_88;
    10'd5:  neuron_6_mul_3_p <= Pix_89;
    10'd6:  neuron_6_mul_3_p <= Pix_90;
    10'd7:  neuron_6_mul_3_p <= Pix_91;
    10'd8:  neuron_6_mul_3_p <= Pix_92;
    10'd9:  neuron_6_mul_3_p <= Pix_93;
    10'd10:  neuron_6_mul_3_p <= Pix_94;
    10'd11:  neuron_6_mul_3_p <= Pix_95;
    10'd12:  neuron_6_mul_3_p <= Pix_96;
    10'd13:  neuron_6_mul_3_p <= Pix_97;
    10'd14:  neuron_6_mul_3_p <= Pix_98;
    10'd15:  neuron_6_mul_3_p <= Pix_99;
    10'd16:  neuron_6_mul_3_p <= Pix_100;
    10'd17:  neuron_6_mul_3_p <= Pix_101;
    10'd18:  neuron_6_mul_3_p <= Pix_102;
    10'd19:  neuron_6_mul_3_p <= Pix_103;
    10'd20:  neuron_6_mul_3_p <= Pix_104;
    10'd21:  neuron_6_mul_3_p <= Pix_105;
    10'd22:  neuron_6_mul_3_p <= Pix_106;
    10'd23:  neuron_6_mul_3_p <= Pix_107;
    10'd24:  neuron_6_mul_3_p <= Pix_108;
    10'd25:  neuron_6_mul_3_p <= Pix_109;
    10'd26:  neuron_6_mul_3_p <= Pix_110;
    10'd27:  neuron_6_mul_3_p <= Pix_111;
    default: neuron_6_mul_3_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_4_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_4_p <= Pix_112;
    10'd1:  neuron_6_mul_4_p <= Pix_113;
    10'd2:  neuron_6_mul_4_p <= Pix_114;
    10'd3:  neuron_6_mul_4_p <= Pix_115;
    10'd4:  neuron_6_mul_4_p <= Pix_116;
    10'd5:  neuron_6_mul_4_p <= Pix_117;
    10'd6:  neuron_6_mul_4_p <= Pix_118;
    10'd7:  neuron_6_mul_4_p <= Pix_119;
    10'd8:  neuron_6_mul_4_p <= Pix_120;
    10'd9:  neuron_6_mul_4_p <= Pix_121;
    10'd10:  neuron_6_mul_4_p <= Pix_122;
    10'd11:  neuron_6_mul_4_p <= Pix_123;
    10'd12:  neuron_6_mul_4_p <= Pix_124;
    10'd13:  neuron_6_mul_4_p <= Pix_125;
    10'd14:  neuron_6_mul_4_p <= Pix_126;
    10'd15:  neuron_6_mul_4_p <= Pix_127;
    10'd16:  neuron_6_mul_4_p <= Pix_128;
    10'd17:  neuron_6_mul_4_p <= Pix_129;
    10'd18:  neuron_6_mul_4_p <= Pix_130;
    10'd19:  neuron_6_mul_4_p <= Pix_131;
    10'd20:  neuron_6_mul_4_p <= Pix_132;
    10'd21:  neuron_6_mul_4_p <= Pix_133;
    10'd22:  neuron_6_mul_4_p <= Pix_134;
    10'd23:  neuron_6_mul_4_p <= Pix_135;
    10'd24:  neuron_6_mul_4_p <= Pix_136;
    10'd25:  neuron_6_mul_4_p <= Pix_137;
    10'd26:  neuron_6_mul_4_p <= Pix_138;
    10'd27:  neuron_6_mul_4_p <= Pix_139;
    default: neuron_6_mul_4_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_5_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_5_p <= Pix_140;
    10'd1:  neuron_6_mul_5_p <= Pix_141;
    10'd2:  neuron_6_mul_5_p <= Pix_142;
    10'd3:  neuron_6_mul_5_p <= Pix_143;
    10'd4:  neuron_6_mul_5_p <= Pix_144;
    10'd5:  neuron_6_mul_5_p <= Pix_145;
    10'd6:  neuron_6_mul_5_p <= Pix_146;
    10'd7:  neuron_6_mul_5_p <= Pix_147;
    10'd8:  neuron_6_mul_5_p <= Pix_148;
    10'd9:  neuron_6_mul_5_p <= Pix_149;
    10'd10:  neuron_6_mul_5_p <= Pix_150;
    10'd11:  neuron_6_mul_5_p <= Pix_151;
    10'd12:  neuron_6_mul_5_p <= Pix_152;
    10'd13:  neuron_6_mul_5_p <= Pix_153;
    10'd14:  neuron_6_mul_5_p <= Pix_154;
    10'd15:  neuron_6_mul_5_p <= Pix_155;
    10'd16:  neuron_6_mul_5_p <= Pix_156;
    10'd17:  neuron_6_mul_5_p <= Pix_157;
    10'd18:  neuron_6_mul_5_p <= Pix_158;
    10'd19:  neuron_6_mul_5_p <= Pix_159;
    10'd20:  neuron_6_mul_5_p <= Pix_160;
    10'd21:  neuron_6_mul_5_p <= Pix_161;
    10'd22:  neuron_6_mul_5_p <= Pix_162;
    10'd23:  neuron_6_mul_5_p <= Pix_163;
    10'd24:  neuron_6_mul_5_p <= Pix_164;
    10'd25:  neuron_6_mul_5_p <= Pix_165;
    10'd26:  neuron_6_mul_5_p <= Pix_166;
    10'd27:  neuron_6_mul_5_p <= Pix_167;
    default: neuron_6_mul_5_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_6_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_6_p <= Pix_168;
    10'd1:  neuron_6_mul_6_p <= Pix_169;
    10'd2:  neuron_6_mul_6_p <= Pix_170;
    10'd3:  neuron_6_mul_6_p <= Pix_171;
    10'd4:  neuron_6_mul_6_p <= Pix_172;
    10'd5:  neuron_6_mul_6_p <= Pix_173;
    10'd6:  neuron_6_mul_6_p <= Pix_174;
    10'd7:  neuron_6_mul_6_p <= Pix_175;
    10'd8:  neuron_6_mul_6_p <= Pix_176;
    10'd9:  neuron_6_mul_6_p <= Pix_177;
    10'd10:  neuron_6_mul_6_p <= Pix_178;
    10'd11:  neuron_6_mul_6_p <= Pix_179;
    10'd12:  neuron_6_mul_6_p <= Pix_180;
    10'd13:  neuron_6_mul_6_p <= Pix_181;
    10'd14:  neuron_6_mul_6_p <= Pix_182;
    10'd15:  neuron_6_mul_6_p <= Pix_183;
    10'd16:  neuron_6_mul_6_p <= Pix_184;
    10'd17:  neuron_6_mul_6_p <= Pix_185;
    10'd18:  neuron_6_mul_6_p <= Pix_186;
    10'd19:  neuron_6_mul_6_p <= Pix_187;
    10'd20:  neuron_6_mul_6_p <= Pix_188;
    10'd21:  neuron_6_mul_6_p <= Pix_189;
    10'd22:  neuron_6_mul_6_p <= Pix_190;
    10'd23:  neuron_6_mul_6_p <= Pix_191;
    10'd24:  neuron_6_mul_6_p <= Pix_192;
    10'd25:  neuron_6_mul_6_p <= Pix_193;
    10'd26:  neuron_6_mul_6_p <= Pix_194;
    10'd27:  neuron_6_mul_6_p <= Pix_195;
    default: neuron_6_mul_6_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_7_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_7_p <= Pix_196;
    10'd1:  neuron_6_mul_7_p <= Pix_197;
    10'd2:  neuron_6_mul_7_p <= Pix_198;
    10'd3:  neuron_6_mul_7_p <= Pix_199;
    10'd4:  neuron_6_mul_7_p <= Pix_200;
    10'd5:  neuron_6_mul_7_p <= Pix_201;
    10'd6:  neuron_6_mul_7_p <= Pix_202;
    10'd7:  neuron_6_mul_7_p <= Pix_203;
    10'd8:  neuron_6_mul_7_p <= Pix_204;
    10'd9:  neuron_6_mul_7_p <= Pix_205;
    10'd10:  neuron_6_mul_7_p <= Pix_206;
    10'd11:  neuron_6_mul_7_p <= Pix_207;
    10'd12:  neuron_6_mul_7_p <= Pix_208;
    10'd13:  neuron_6_mul_7_p <= Pix_209;
    10'd14:  neuron_6_mul_7_p <= Pix_210;
    10'd15:  neuron_6_mul_7_p <= Pix_211;
    10'd16:  neuron_6_mul_7_p <= Pix_212;
    10'd17:  neuron_6_mul_7_p <= Pix_213;
    10'd18:  neuron_6_mul_7_p <= Pix_214;
    10'd19:  neuron_6_mul_7_p <= Pix_215;
    10'd20:  neuron_6_mul_7_p <= Pix_216;
    10'd21:  neuron_6_mul_7_p <= Pix_217;
    10'd22:  neuron_6_mul_7_p <= Pix_218;
    10'd23:  neuron_6_mul_7_p <= Pix_219;
    10'd24:  neuron_6_mul_7_p <= Pix_220;
    10'd25:  neuron_6_mul_7_p <= Pix_221;
    10'd26:  neuron_6_mul_7_p <= Pix_222;
    10'd27:  neuron_6_mul_7_p <= Pix_223;
    default: neuron_6_mul_7_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_8_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_8_p <= Pix_224;
    10'd1:  neuron_6_mul_8_p <= Pix_225;
    10'd2:  neuron_6_mul_8_p <= Pix_226;
    10'd3:  neuron_6_mul_8_p <= Pix_227;
    10'd4:  neuron_6_mul_8_p <= Pix_228;
    10'd5:  neuron_6_mul_8_p <= Pix_229;
    10'd6:  neuron_6_mul_8_p <= Pix_230;
    10'd7:  neuron_6_mul_8_p <= Pix_231;
    10'd8:  neuron_6_mul_8_p <= Pix_232;
    10'd9:  neuron_6_mul_8_p <= Pix_233;
    10'd10:  neuron_6_mul_8_p <= Pix_234;
    10'd11:  neuron_6_mul_8_p <= Pix_235;
    10'd12:  neuron_6_mul_8_p <= Pix_236;
    10'd13:  neuron_6_mul_8_p <= Pix_237;
    10'd14:  neuron_6_mul_8_p <= Pix_238;
    10'd15:  neuron_6_mul_8_p <= Pix_239;
    10'd16:  neuron_6_mul_8_p <= Pix_240;
    10'd17:  neuron_6_mul_8_p <= Pix_241;
    10'd18:  neuron_6_mul_8_p <= Pix_242;
    10'd19:  neuron_6_mul_8_p <= Pix_243;
    10'd20:  neuron_6_mul_8_p <= Pix_244;
    10'd21:  neuron_6_mul_8_p <= Pix_245;
    10'd22:  neuron_6_mul_8_p <= Pix_246;
    10'd23:  neuron_6_mul_8_p <= Pix_247;
    10'd24:  neuron_6_mul_8_p <= Pix_248;
    10'd25:  neuron_6_mul_8_p <= Pix_249;
    10'd26:  neuron_6_mul_8_p <= Pix_250;
    10'd27:  neuron_6_mul_8_p <= Pix_251;
    default: neuron_6_mul_8_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_9_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_9_p <= Pix_252;
    10'd1:  neuron_6_mul_9_p <= Pix_253;
    10'd2:  neuron_6_mul_9_p <= Pix_254;
    10'd3:  neuron_6_mul_9_p <= Pix_255;
    10'd4:  neuron_6_mul_9_p <= Pix_256;
    10'd5:  neuron_6_mul_9_p <= Pix_257;
    10'd6:  neuron_6_mul_9_p <= Pix_258;
    10'd7:  neuron_6_mul_9_p <= Pix_259;
    10'd8:  neuron_6_mul_9_p <= Pix_260;
    10'd9:  neuron_6_mul_9_p <= Pix_261;
    10'd10:  neuron_6_mul_9_p <= Pix_262;
    10'd11:  neuron_6_mul_9_p <= Pix_263;
    10'd12:  neuron_6_mul_9_p <= Pix_264;
    10'd13:  neuron_6_mul_9_p <= Pix_265;
    10'd14:  neuron_6_mul_9_p <= Pix_266;
    10'd15:  neuron_6_mul_9_p <= Pix_267;
    10'd16:  neuron_6_mul_9_p <= Pix_268;
    10'd17:  neuron_6_mul_9_p <= Pix_269;
    10'd18:  neuron_6_mul_9_p <= Pix_270;
    10'd19:  neuron_6_mul_9_p <= Pix_271;
    10'd20:  neuron_6_mul_9_p <= Pix_272;
    10'd21:  neuron_6_mul_9_p <= Pix_273;
    10'd22:  neuron_6_mul_9_p <= Pix_274;
    10'd23:  neuron_6_mul_9_p <= Pix_275;
    10'd24:  neuron_6_mul_9_p <= Pix_276;
    10'd25:  neuron_6_mul_9_p <= Pix_277;
    10'd26:  neuron_6_mul_9_p <= Pix_278;
    10'd27:  neuron_6_mul_9_p <= Pix_279;
    default: neuron_6_mul_9_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_10_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_10_p <= Pix_280;
    10'd1:  neuron_6_mul_10_p <= Pix_281;
    10'd2:  neuron_6_mul_10_p <= Pix_282;
    10'd3:  neuron_6_mul_10_p <= Pix_283;
    10'd4:  neuron_6_mul_10_p <= Pix_284;
    10'd5:  neuron_6_mul_10_p <= Pix_285;
    10'd6:  neuron_6_mul_10_p <= Pix_286;
    10'd7:  neuron_6_mul_10_p <= Pix_287;
    10'd8:  neuron_6_mul_10_p <= Pix_288;
    10'd9:  neuron_6_mul_10_p <= Pix_289;
    10'd10:  neuron_6_mul_10_p <= Pix_290;
    10'd11:  neuron_6_mul_10_p <= Pix_291;
    10'd12:  neuron_6_mul_10_p <= Pix_292;
    10'd13:  neuron_6_mul_10_p <= Pix_293;
    10'd14:  neuron_6_mul_10_p <= Pix_294;
    10'd15:  neuron_6_mul_10_p <= Pix_295;
    10'd16:  neuron_6_mul_10_p <= Pix_296;
    10'd17:  neuron_6_mul_10_p <= Pix_297;
    10'd18:  neuron_6_mul_10_p <= Pix_298;
    10'd19:  neuron_6_mul_10_p <= Pix_299;
    10'd20:  neuron_6_mul_10_p <= Pix_300;
    10'd21:  neuron_6_mul_10_p <= Pix_301;
    10'd22:  neuron_6_mul_10_p <= Pix_302;
    10'd23:  neuron_6_mul_10_p <= Pix_303;
    10'd24:  neuron_6_mul_10_p <= Pix_304;
    10'd25:  neuron_6_mul_10_p <= Pix_305;
    10'd26:  neuron_6_mul_10_p <= Pix_306;
    10'd27:  neuron_6_mul_10_p <= Pix_307;
    default: neuron_6_mul_10_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_11_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_11_p <= Pix_308;
    10'd1:  neuron_6_mul_11_p <= Pix_309;
    10'd2:  neuron_6_mul_11_p <= Pix_310;
    10'd3:  neuron_6_mul_11_p <= Pix_311;
    10'd4:  neuron_6_mul_11_p <= Pix_312;
    10'd5:  neuron_6_mul_11_p <= Pix_313;
    10'd6:  neuron_6_mul_11_p <= Pix_314;
    10'd7:  neuron_6_mul_11_p <= Pix_315;
    10'd8:  neuron_6_mul_11_p <= Pix_316;
    10'd9:  neuron_6_mul_11_p <= Pix_317;
    10'd10:  neuron_6_mul_11_p <= Pix_318;
    10'd11:  neuron_6_mul_11_p <= Pix_319;
    10'd12:  neuron_6_mul_11_p <= Pix_320;
    10'd13:  neuron_6_mul_11_p <= Pix_321;
    10'd14:  neuron_6_mul_11_p <= Pix_322;
    10'd15:  neuron_6_mul_11_p <= Pix_323;
    10'd16:  neuron_6_mul_11_p <= Pix_324;
    10'd17:  neuron_6_mul_11_p <= Pix_325;
    10'd18:  neuron_6_mul_11_p <= Pix_326;
    10'd19:  neuron_6_mul_11_p <= Pix_327;
    10'd20:  neuron_6_mul_11_p <= Pix_328;
    10'd21:  neuron_6_mul_11_p <= Pix_329;
    10'd22:  neuron_6_mul_11_p <= Pix_330;
    10'd23:  neuron_6_mul_11_p <= Pix_331;
    10'd24:  neuron_6_mul_11_p <= Pix_332;
    10'd25:  neuron_6_mul_11_p <= Pix_333;
    10'd26:  neuron_6_mul_11_p <= Pix_334;
    10'd27:  neuron_6_mul_11_p <= Pix_335;
    default: neuron_6_mul_11_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_12_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_12_p <= Pix_336;
    10'd1:  neuron_6_mul_12_p <= Pix_337;
    10'd2:  neuron_6_mul_12_p <= Pix_338;
    10'd3:  neuron_6_mul_12_p <= Pix_339;
    10'd4:  neuron_6_mul_12_p <= Pix_340;
    10'd5:  neuron_6_mul_12_p <= Pix_341;
    10'd6:  neuron_6_mul_12_p <= Pix_342;
    10'd7:  neuron_6_mul_12_p <= Pix_343;
    10'd8:  neuron_6_mul_12_p <= Pix_344;
    10'd9:  neuron_6_mul_12_p <= Pix_345;
    10'd10:  neuron_6_mul_12_p <= Pix_346;
    10'd11:  neuron_6_mul_12_p <= Pix_347;
    10'd12:  neuron_6_mul_12_p <= Pix_348;
    10'd13:  neuron_6_mul_12_p <= Pix_349;
    10'd14:  neuron_6_mul_12_p <= Pix_350;
    10'd15:  neuron_6_mul_12_p <= Pix_351;
    10'd16:  neuron_6_mul_12_p <= Pix_352;
    10'd17:  neuron_6_mul_12_p <= Pix_353;
    10'd18:  neuron_6_mul_12_p <= Pix_354;
    10'd19:  neuron_6_mul_12_p <= Pix_355;
    10'd20:  neuron_6_mul_12_p <= Pix_356;
    10'd21:  neuron_6_mul_12_p <= Pix_357;
    10'd22:  neuron_6_mul_12_p <= Pix_358;
    10'd23:  neuron_6_mul_12_p <= Pix_359;
    10'd24:  neuron_6_mul_12_p <= Pix_360;
    10'd25:  neuron_6_mul_12_p <= Pix_361;
    10'd26:  neuron_6_mul_12_p <= Pix_362;
    10'd27:  neuron_6_mul_12_p <= Pix_363;
    default: neuron_6_mul_12_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_13_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_13_p <= Pix_364;
    10'd1:  neuron_6_mul_13_p <= Pix_365;
    10'd2:  neuron_6_mul_13_p <= Pix_366;
    10'd3:  neuron_6_mul_13_p <= Pix_367;
    10'd4:  neuron_6_mul_13_p <= Pix_368;
    10'd5:  neuron_6_mul_13_p <= Pix_369;
    10'd6:  neuron_6_mul_13_p <= Pix_370;
    10'd7:  neuron_6_mul_13_p <= Pix_371;
    10'd8:  neuron_6_mul_13_p <= Pix_372;
    10'd9:  neuron_6_mul_13_p <= Pix_373;
    10'd10:  neuron_6_mul_13_p <= Pix_374;
    10'd11:  neuron_6_mul_13_p <= Pix_375;
    10'd12:  neuron_6_mul_13_p <= Pix_376;
    10'd13:  neuron_6_mul_13_p <= Pix_377;
    10'd14:  neuron_6_mul_13_p <= Pix_378;
    10'd15:  neuron_6_mul_13_p <= Pix_379;
    10'd16:  neuron_6_mul_13_p <= Pix_380;
    10'd17:  neuron_6_mul_13_p <= Pix_381;
    10'd18:  neuron_6_mul_13_p <= Pix_382;
    10'd19:  neuron_6_mul_13_p <= Pix_383;
    10'd20:  neuron_6_mul_13_p <= Pix_384;
    10'd21:  neuron_6_mul_13_p <= Pix_385;
    10'd22:  neuron_6_mul_13_p <= Pix_386;
    10'd23:  neuron_6_mul_13_p <= Pix_387;
    10'd24:  neuron_6_mul_13_p <= Pix_388;
    10'd25:  neuron_6_mul_13_p <= Pix_389;
    10'd26:  neuron_6_mul_13_p <= Pix_390;
    10'd27:  neuron_6_mul_13_p <= Pix_391;
    default: neuron_6_mul_13_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_14_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_14_p <= Pix_392;
    10'd1:  neuron_6_mul_14_p <= Pix_393;
    10'd2:  neuron_6_mul_14_p <= Pix_394;
    10'd3:  neuron_6_mul_14_p <= Pix_395;
    10'd4:  neuron_6_mul_14_p <= Pix_396;
    10'd5:  neuron_6_mul_14_p <= Pix_397;
    10'd6:  neuron_6_mul_14_p <= Pix_398;
    10'd7:  neuron_6_mul_14_p <= Pix_399;
    10'd8:  neuron_6_mul_14_p <= Pix_400;
    10'd9:  neuron_6_mul_14_p <= Pix_401;
    10'd10:  neuron_6_mul_14_p <= Pix_402;
    10'd11:  neuron_6_mul_14_p <= Pix_403;
    10'd12:  neuron_6_mul_14_p <= Pix_404;
    10'd13:  neuron_6_mul_14_p <= Pix_405;
    10'd14:  neuron_6_mul_14_p <= Pix_406;
    10'd15:  neuron_6_mul_14_p <= Pix_407;
    10'd16:  neuron_6_mul_14_p <= Pix_408;
    10'd17:  neuron_6_mul_14_p <= Pix_409;
    10'd18:  neuron_6_mul_14_p <= Pix_410;
    10'd19:  neuron_6_mul_14_p <= Pix_411;
    10'd20:  neuron_6_mul_14_p <= Pix_412;
    10'd21:  neuron_6_mul_14_p <= Pix_413;
    10'd22:  neuron_6_mul_14_p <= Pix_414;
    10'd23:  neuron_6_mul_14_p <= Pix_415;
    10'd24:  neuron_6_mul_14_p <= Pix_416;
    10'd25:  neuron_6_mul_14_p <= Pix_417;
    10'd26:  neuron_6_mul_14_p <= Pix_418;
    10'd27:  neuron_6_mul_14_p <= Pix_419;
    default: neuron_6_mul_14_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_15_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_15_p <= Pix_420;
    10'd1:  neuron_6_mul_15_p <= Pix_421;
    10'd2:  neuron_6_mul_15_p <= Pix_422;
    10'd3:  neuron_6_mul_15_p <= Pix_423;
    10'd4:  neuron_6_mul_15_p <= Pix_424;
    10'd5:  neuron_6_mul_15_p <= Pix_425;
    10'd6:  neuron_6_mul_15_p <= Pix_426;
    10'd7:  neuron_6_mul_15_p <= Pix_427;
    10'd8:  neuron_6_mul_15_p <= Pix_428;
    10'd9:  neuron_6_mul_15_p <= Pix_429;
    10'd10:  neuron_6_mul_15_p <= Pix_430;
    10'd11:  neuron_6_mul_15_p <= Pix_431;
    10'd12:  neuron_6_mul_15_p <= Pix_432;
    10'd13:  neuron_6_mul_15_p <= Pix_433;
    10'd14:  neuron_6_mul_15_p <= Pix_434;
    10'd15:  neuron_6_mul_15_p <= Pix_435;
    10'd16:  neuron_6_mul_15_p <= Pix_436;
    10'd17:  neuron_6_mul_15_p <= Pix_437;
    10'd18:  neuron_6_mul_15_p <= Pix_438;
    10'd19:  neuron_6_mul_15_p <= Pix_439;
    10'd20:  neuron_6_mul_15_p <= Pix_440;
    10'd21:  neuron_6_mul_15_p <= Pix_441;
    10'd22:  neuron_6_mul_15_p <= Pix_442;
    10'd23:  neuron_6_mul_15_p <= Pix_443;
    10'd24:  neuron_6_mul_15_p <= Pix_444;
    10'd25:  neuron_6_mul_15_p <= Pix_445;
    10'd26:  neuron_6_mul_15_p <= Pix_446;
    10'd27:  neuron_6_mul_15_p <= Pix_447;
    default: neuron_6_mul_15_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_16_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_16_p <= Pix_448;
    10'd1:  neuron_6_mul_16_p <= Pix_449;
    10'd2:  neuron_6_mul_16_p <= Pix_450;
    10'd3:  neuron_6_mul_16_p <= Pix_451;
    10'd4:  neuron_6_mul_16_p <= Pix_452;
    10'd5:  neuron_6_mul_16_p <= Pix_453;
    10'd6:  neuron_6_mul_16_p <= Pix_454;
    10'd7:  neuron_6_mul_16_p <= Pix_455;
    10'd8:  neuron_6_mul_16_p <= Pix_456;
    10'd9:  neuron_6_mul_16_p <= Pix_457;
    10'd10:  neuron_6_mul_16_p <= Pix_458;
    10'd11:  neuron_6_mul_16_p <= Pix_459;
    10'd12:  neuron_6_mul_16_p <= Pix_460;
    10'd13:  neuron_6_mul_16_p <= Pix_461;
    10'd14:  neuron_6_mul_16_p <= Pix_462;
    10'd15:  neuron_6_mul_16_p <= Pix_463;
    10'd16:  neuron_6_mul_16_p <= Pix_464;
    10'd17:  neuron_6_mul_16_p <= Pix_465;
    10'd18:  neuron_6_mul_16_p <= Pix_466;
    10'd19:  neuron_6_mul_16_p <= Pix_467;
    10'd20:  neuron_6_mul_16_p <= Pix_468;
    10'd21:  neuron_6_mul_16_p <= Pix_469;
    10'd22:  neuron_6_mul_16_p <= Pix_470;
    10'd23:  neuron_6_mul_16_p <= Pix_471;
    10'd24:  neuron_6_mul_16_p <= Pix_472;
    10'd25:  neuron_6_mul_16_p <= Pix_473;
    10'd26:  neuron_6_mul_16_p <= Pix_474;
    10'd27:  neuron_6_mul_16_p <= Pix_475;
    default: neuron_6_mul_16_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_17_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_17_p <= Pix_476;
    10'd1:  neuron_6_mul_17_p <= Pix_477;
    10'd2:  neuron_6_mul_17_p <= Pix_478;
    10'd3:  neuron_6_mul_17_p <= Pix_479;
    10'd4:  neuron_6_mul_17_p <= Pix_480;
    10'd5:  neuron_6_mul_17_p <= Pix_481;
    10'd6:  neuron_6_mul_17_p <= Pix_482;
    10'd7:  neuron_6_mul_17_p <= Pix_483;
    10'd8:  neuron_6_mul_17_p <= Pix_484;
    10'd9:  neuron_6_mul_17_p <= Pix_485;
    10'd10:  neuron_6_mul_17_p <= Pix_486;
    10'd11:  neuron_6_mul_17_p <= Pix_487;
    10'd12:  neuron_6_mul_17_p <= Pix_488;
    10'd13:  neuron_6_mul_17_p <= Pix_489;
    10'd14:  neuron_6_mul_17_p <= Pix_490;
    10'd15:  neuron_6_mul_17_p <= Pix_491;
    10'd16:  neuron_6_mul_17_p <= Pix_492;
    10'd17:  neuron_6_mul_17_p <= Pix_493;
    10'd18:  neuron_6_mul_17_p <= Pix_494;
    10'd19:  neuron_6_mul_17_p <= Pix_495;
    10'd20:  neuron_6_mul_17_p <= Pix_496;
    10'd21:  neuron_6_mul_17_p <= Pix_497;
    10'd22:  neuron_6_mul_17_p <= Pix_498;
    10'd23:  neuron_6_mul_17_p <= Pix_499;
    10'd24:  neuron_6_mul_17_p <= Pix_500;
    10'd25:  neuron_6_mul_17_p <= Pix_501;
    10'd26:  neuron_6_mul_17_p <= Pix_502;
    10'd27:  neuron_6_mul_17_p <= Pix_503;
    default: neuron_6_mul_17_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_18_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_18_p <= Pix_504;
    10'd1:  neuron_6_mul_18_p <= Pix_505;
    10'd2:  neuron_6_mul_18_p <= Pix_506;
    10'd3:  neuron_6_mul_18_p <= Pix_507;
    10'd4:  neuron_6_mul_18_p <= Pix_508;
    10'd5:  neuron_6_mul_18_p <= Pix_509;
    10'd6:  neuron_6_mul_18_p <= Pix_510;
    10'd7:  neuron_6_mul_18_p <= Pix_511;
    10'd8:  neuron_6_mul_18_p <= Pix_512;
    10'd9:  neuron_6_mul_18_p <= Pix_513;
    10'd10:  neuron_6_mul_18_p <= Pix_514;
    10'd11:  neuron_6_mul_18_p <= Pix_515;
    10'd12:  neuron_6_mul_18_p <= Pix_516;
    10'd13:  neuron_6_mul_18_p <= Pix_517;
    10'd14:  neuron_6_mul_18_p <= Pix_518;
    10'd15:  neuron_6_mul_18_p <= Pix_519;
    10'd16:  neuron_6_mul_18_p <= Pix_520;
    10'd17:  neuron_6_mul_18_p <= Pix_521;
    10'd18:  neuron_6_mul_18_p <= Pix_522;
    10'd19:  neuron_6_mul_18_p <= Pix_523;
    10'd20:  neuron_6_mul_18_p <= Pix_524;
    10'd21:  neuron_6_mul_18_p <= Pix_525;
    10'd22:  neuron_6_mul_18_p <= Pix_526;
    10'd23:  neuron_6_mul_18_p <= Pix_527;
    10'd24:  neuron_6_mul_18_p <= Pix_528;
    10'd25:  neuron_6_mul_18_p <= Pix_529;
    10'd26:  neuron_6_mul_18_p <= Pix_530;
    10'd27:  neuron_6_mul_18_p <= Pix_531;
    default: neuron_6_mul_18_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_19_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_19_p <= Pix_532;
    10'd1:  neuron_6_mul_19_p <= Pix_533;
    10'd2:  neuron_6_mul_19_p <= Pix_534;
    10'd3:  neuron_6_mul_19_p <= Pix_535;
    10'd4:  neuron_6_mul_19_p <= Pix_536;
    10'd5:  neuron_6_mul_19_p <= Pix_537;
    10'd6:  neuron_6_mul_19_p <= Pix_538;
    10'd7:  neuron_6_mul_19_p <= Pix_539;
    10'd8:  neuron_6_mul_19_p <= Pix_540;
    10'd9:  neuron_6_mul_19_p <= Pix_541;
    10'd10:  neuron_6_mul_19_p <= Pix_542;
    10'd11:  neuron_6_mul_19_p <= Pix_543;
    10'd12:  neuron_6_mul_19_p <= Pix_544;
    10'd13:  neuron_6_mul_19_p <= Pix_545;
    10'd14:  neuron_6_mul_19_p <= Pix_546;
    10'd15:  neuron_6_mul_19_p <= Pix_547;
    10'd16:  neuron_6_mul_19_p <= Pix_548;
    10'd17:  neuron_6_mul_19_p <= Pix_549;
    10'd18:  neuron_6_mul_19_p <= Pix_550;
    10'd19:  neuron_6_mul_19_p <= Pix_551;
    10'd20:  neuron_6_mul_19_p <= Pix_552;
    10'd21:  neuron_6_mul_19_p <= Pix_553;
    10'd22:  neuron_6_mul_19_p <= Pix_554;
    10'd23:  neuron_6_mul_19_p <= Pix_555;
    10'd24:  neuron_6_mul_19_p <= Pix_556;
    10'd25:  neuron_6_mul_19_p <= Pix_557;
    10'd26:  neuron_6_mul_19_p <= Pix_558;
    10'd27:  neuron_6_mul_19_p <= Pix_559;
    default: neuron_6_mul_19_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_20_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_20_p <= Pix_560;
    10'd1:  neuron_6_mul_20_p <= Pix_561;
    10'd2:  neuron_6_mul_20_p <= Pix_562;
    10'd3:  neuron_6_mul_20_p <= Pix_563;
    10'd4:  neuron_6_mul_20_p <= Pix_564;
    10'd5:  neuron_6_mul_20_p <= Pix_565;
    10'd6:  neuron_6_mul_20_p <= Pix_566;
    10'd7:  neuron_6_mul_20_p <= Pix_567;
    10'd8:  neuron_6_mul_20_p <= Pix_568;
    10'd9:  neuron_6_mul_20_p <= Pix_569;
    10'd10:  neuron_6_mul_20_p <= Pix_570;
    10'd11:  neuron_6_mul_20_p <= Pix_571;
    10'd12:  neuron_6_mul_20_p <= Pix_572;
    10'd13:  neuron_6_mul_20_p <= Pix_573;
    10'd14:  neuron_6_mul_20_p <= Pix_574;
    10'd15:  neuron_6_mul_20_p <= Pix_575;
    10'd16:  neuron_6_mul_20_p <= Pix_576;
    10'd17:  neuron_6_mul_20_p <= Pix_577;
    10'd18:  neuron_6_mul_20_p <= Pix_578;
    10'd19:  neuron_6_mul_20_p <= Pix_579;
    10'd20:  neuron_6_mul_20_p <= Pix_580;
    10'd21:  neuron_6_mul_20_p <= Pix_581;
    10'd22:  neuron_6_mul_20_p <= Pix_582;
    10'd23:  neuron_6_mul_20_p <= Pix_583;
    10'd24:  neuron_6_mul_20_p <= Pix_584;
    10'd25:  neuron_6_mul_20_p <= Pix_585;
    10'd26:  neuron_6_mul_20_p <= Pix_586;
    10'd27:  neuron_6_mul_20_p <= Pix_587;
    default: neuron_6_mul_20_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_21_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_21_p <= Pix_588;
    10'd1:  neuron_6_mul_21_p <= Pix_589;
    10'd2:  neuron_6_mul_21_p <= Pix_590;
    10'd3:  neuron_6_mul_21_p <= Pix_591;
    10'd4:  neuron_6_mul_21_p <= Pix_592;
    10'd5:  neuron_6_mul_21_p <= Pix_593;
    10'd6:  neuron_6_mul_21_p <= Pix_594;
    10'd7:  neuron_6_mul_21_p <= Pix_595;
    10'd8:  neuron_6_mul_21_p <= Pix_596;
    10'd9:  neuron_6_mul_21_p <= Pix_597;
    10'd10:  neuron_6_mul_21_p <= Pix_598;
    10'd11:  neuron_6_mul_21_p <= Pix_599;
    10'd12:  neuron_6_mul_21_p <= Pix_600;
    10'd13:  neuron_6_mul_21_p <= Pix_601;
    10'd14:  neuron_6_mul_21_p <= Pix_602;
    10'd15:  neuron_6_mul_21_p <= Pix_603;
    10'd16:  neuron_6_mul_21_p <= Pix_604;
    10'd17:  neuron_6_mul_21_p <= Pix_605;
    10'd18:  neuron_6_mul_21_p <= Pix_606;
    10'd19:  neuron_6_mul_21_p <= Pix_607;
    10'd20:  neuron_6_mul_21_p <= Pix_608;
    10'd21:  neuron_6_mul_21_p <= Pix_609;
    10'd22:  neuron_6_mul_21_p <= Pix_610;
    10'd23:  neuron_6_mul_21_p <= Pix_611;
    10'd24:  neuron_6_mul_21_p <= Pix_612;
    10'd25:  neuron_6_mul_21_p <= Pix_613;
    10'd26:  neuron_6_mul_21_p <= Pix_614;
    10'd27:  neuron_6_mul_21_p <= Pix_615;
    default: neuron_6_mul_21_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_22_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_22_p <= Pix_616;
    10'd1:  neuron_6_mul_22_p <= Pix_617;
    10'd2:  neuron_6_mul_22_p <= Pix_618;
    10'd3:  neuron_6_mul_22_p <= Pix_619;
    10'd4:  neuron_6_mul_22_p <= Pix_620;
    10'd5:  neuron_6_mul_22_p <= Pix_621;
    10'd6:  neuron_6_mul_22_p <= Pix_622;
    10'd7:  neuron_6_mul_22_p <= Pix_623;
    10'd8:  neuron_6_mul_22_p <= Pix_624;
    10'd9:  neuron_6_mul_22_p <= Pix_625;
    10'd10:  neuron_6_mul_22_p <= Pix_626;
    10'd11:  neuron_6_mul_22_p <= Pix_627;
    10'd12:  neuron_6_mul_22_p <= Pix_628;
    10'd13:  neuron_6_mul_22_p <= Pix_629;
    10'd14:  neuron_6_mul_22_p <= Pix_630;
    10'd15:  neuron_6_mul_22_p <= Pix_631;
    10'd16:  neuron_6_mul_22_p <= Pix_632;
    10'd17:  neuron_6_mul_22_p <= Pix_633;
    10'd18:  neuron_6_mul_22_p <= Pix_634;
    10'd19:  neuron_6_mul_22_p <= Pix_635;
    10'd20:  neuron_6_mul_22_p <= Pix_636;
    10'd21:  neuron_6_mul_22_p <= Pix_637;
    10'd22:  neuron_6_mul_22_p <= Pix_638;
    10'd23:  neuron_6_mul_22_p <= Pix_639;
    10'd24:  neuron_6_mul_22_p <= Pix_640;
    10'd25:  neuron_6_mul_22_p <= Pix_641;
    10'd26:  neuron_6_mul_22_p <= Pix_642;
    10'd27:  neuron_6_mul_22_p <= Pix_643;
    default: neuron_6_mul_22_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_23_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_23_p <= Pix_644;
    10'd1:  neuron_6_mul_23_p <= Pix_645;
    10'd2:  neuron_6_mul_23_p <= Pix_646;
    10'd3:  neuron_6_mul_23_p <= Pix_647;
    10'd4:  neuron_6_mul_23_p <= Pix_648;
    10'd5:  neuron_6_mul_23_p <= Pix_649;
    10'd6:  neuron_6_mul_23_p <= Pix_650;
    10'd7:  neuron_6_mul_23_p <= Pix_651;
    10'd8:  neuron_6_mul_23_p <= Pix_652;
    10'd9:  neuron_6_mul_23_p <= Pix_653;
    10'd10:  neuron_6_mul_23_p <= Pix_654;
    10'd11:  neuron_6_mul_23_p <= Pix_655;
    10'd12:  neuron_6_mul_23_p <= Pix_656;
    10'd13:  neuron_6_mul_23_p <= Pix_657;
    10'd14:  neuron_6_mul_23_p <= Pix_658;
    10'd15:  neuron_6_mul_23_p <= Pix_659;
    10'd16:  neuron_6_mul_23_p <= Pix_660;
    10'd17:  neuron_6_mul_23_p <= Pix_661;
    10'd18:  neuron_6_mul_23_p <= Pix_662;
    10'd19:  neuron_6_mul_23_p <= Pix_663;
    10'd20:  neuron_6_mul_23_p <= Pix_664;
    10'd21:  neuron_6_mul_23_p <= Pix_665;
    10'd22:  neuron_6_mul_23_p <= Pix_666;
    10'd23:  neuron_6_mul_23_p <= Pix_667;
    10'd24:  neuron_6_mul_23_p <= Pix_668;
    10'd25:  neuron_6_mul_23_p <= Pix_669;
    10'd26:  neuron_6_mul_23_p <= Pix_670;
    10'd27:  neuron_6_mul_23_p <= Pix_671;
    default: neuron_6_mul_23_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_24_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_24_p <= Pix_672;
    10'd1:  neuron_6_mul_24_p <= Pix_673;
    10'd2:  neuron_6_mul_24_p <= Pix_674;
    10'd3:  neuron_6_mul_24_p <= Pix_675;
    10'd4:  neuron_6_mul_24_p <= Pix_676;
    10'd5:  neuron_6_mul_24_p <= Pix_677;
    10'd6:  neuron_6_mul_24_p <= Pix_678;
    10'd7:  neuron_6_mul_24_p <= Pix_679;
    10'd8:  neuron_6_mul_24_p <= Pix_680;
    10'd9:  neuron_6_mul_24_p <= Pix_681;
    10'd10:  neuron_6_mul_24_p <= Pix_682;
    10'd11:  neuron_6_mul_24_p <= Pix_683;
    10'd12:  neuron_6_mul_24_p <= Pix_684;
    10'd13:  neuron_6_mul_24_p <= Pix_685;
    10'd14:  neuron_6_mul_24_p <= Pix_686;
    10'd15:  neuron_6_mul_24_p <= Pix_687;
    10'd16:  neuron_6_mul_24_p <= Pix_688;
    10'd17:  neuron_6_mul_24_p <= Pix_689;
    10'd18:  neuron_6_mul_24_p <= Pix_690;
    10'd19:  neuron_6_mul_24_p <= Pix_691;
    10'd20:  neuron_6_mul_24_p <= Pix_692;
    10'd21:  neuron_6_mul_24_p <= Pix_693;
    10'd22:  neuron_6_mul_24_p <= Pix_694;
    10'd23:  neuron_6_mul_24_p <= Pix_695;
    10'd24:  neuron_6_mul_24_p <= Pix_696;
    10'd25:  neuron_6_mul_24_p <= Pix_697;
    10'd26:  neuron_6_mul_24_p <= Pix_698;
    10'd27:  neuron_6_mul_24_p <= Pix_699;
    default: neuron_6_mul_24_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_25_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_25_p <= Pix_700;
    10'd1:  neuron_6_mul_25_p <= Pix_701;
    10'd2:  neuron_6_mul_25_p <= Pix_702;
    10'd3:  neuron_6_mul_25_p <= Pix_703;
    10'd4:  neuron_6_mul_25_p <= Pix_704;
    10'd5:  neuron_6_mul_25_p <= Pix_705;
    10'd6:  neuron_6_mul_25_p <= Pix_706;
    10'd7:  neuron_6_mul_25_p <= Pix_707;
    10'd8:  neuron_6_mul_25_p <= Pix_708;
    10'd9:  neuron_6_mul_25_p <= Pix_709;
    10'd10:  neuron_6_mul_25_p <= Pix_710;
    10'd11:  neuron_6_mul_25_p <= Pix_711;
    10'd12:  neuron_6_mul_25_p <= Pix_712;
    10'd13:  neuron_6_mul_25_p <= Pix_713;
    10'd14:  neuron_6_mul_25_p <= Pix_714;
    10'd15:  neuron_6_mul_25_p <= Pix_715;
    10'd16:  neuron_6_mul_25_p <= Pix_716;
    10'd17:  neuron_6_mul_25_p <= Pix_717;
    10'd18:  neuron_6_mul_25_p <= Pix_718;
    10'd19:  neuron_6_mul_25_p <= Pix_719;
    10'd20:  neuron_6_mul_25_p <= Pix_720;
    10'd21:  neuron_6_mul_25_p <= Pix_721;
    10'd22:  neuron_6_mul_25_p <= Pix_722;
    10'd23:  neuron_6_mul_25_p <= Pix_723;
    10'd24:  neuron_6_mul_25_p <= Pix_724;
    10'd25:  neuron_6_mul_25_p <= Pix_725;
    10'd26:  neuron_6_mul_25_p <= Pix_726;
    10'd27:  neuron_6_mul_25_p <= Pix_727;
    default: neuron_6_mul_25_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_26_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_26_p <= Pix_728;
    10'd1:  neuron_6_mul_26_p <= Pix_729;
    10'd2:  neuron_6_mul_26_p <= Pix_730;
    10'd3:  neuron_6_mul_26_p <= Pix_731;
    10'd4:  neuron_6_mul_26_p <= Pix_732;
    10'd5:  neuron_6_mul_26_p <= Pix_733;
    10'd6:  neuron_6_mul_26_p <= Pix_734;
    10'd7:  neuron_6_mul_26_p <= Pix_735;
    10'd8:  neuron_6_mul_26_p <= Pix_736;
    10'd9:  neuron_6_mul_26_p <= Pix_737;
    10'd10:  neuron_6_mul_26_p <= Pix_738;
    10'd11:  neuron_6_mul_26_p <= Pix_739;
    10'd12:  neuron_6_mul_26_p <= Pix_740;
    10'd13:  neuron_6_mul_26_p <= Pix_741;
    10'd14:  neuron_6_mul_26_p <= Pix_742;
    10'd15:  neuron_6_mul_26_p <= Pix_743;
    10'd16:  neuron_6_mul_26_p <= Pix_744;
    10'd17:  neuron_6_mul_26_p <= Pix_745;
    10'd18:  neuron_6_mul_26_p <= Pix_746;
    10'd19:  neuron_6_mul_26_p <= Pix_747;
    10'd20:  neuron_6_mul_26_p <= Pix_748;
    10'd21:  neuron_6_mul_26_p <= Pix_749;
    10'd22:  neuron_6_mul_26_p <= Pix_750;
    10'd23:  neuron_6_mul_26_p <= Pix_751;
    10'd24:  neuron_6_mul_26_p <= Pix_752;
    10'd25:  neuron_6_mul_26_p <= Pix_753;
    10'd26:  neuron_6_mul_26_p <= Pix_754;
    10'd27:  neuron_6_mul_26_p <= Pix_755;
    default: neuron_6_mul_26_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_6_mul_27_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_6_mul_27_p <= Pix_756;
    10'd1:  neuron_6_mul_27_p <= Pix_757;
    10'd2:  neuron_6_mul_27_p <= Pix_758;
    10'd3:  neuron_6_mul_27_p <= Pix_759;
    10'd4:  neuron_6_mul_27_p <= Pix_760;
    10'd5:  neuron_6_mul_27_p <= Pix_761;
    10'd6:  neuron_6_mul_27_p <= Pix_762;
    10'd7:  neuron_6_mul_27_p <= Pix_763;
    10'd8:  neuron_6_mul_27_p <= Pix_764;
    10'd9:  neuron_6_mul_27_p <= Pix_765;
    10'd10:  neuron_6_mul_27_p <= Pix_766;
    10'd11:  neuron_6_mul_27_p <= Pix_767;
    10'd12:  neuron_6_mul_27_p <= Pix_768;
    10'd13:  neuron_6_mul_27_p <= Pix_769;
    10'd14:  neuron_6_mul_27_p <= Pix_770;
    10'd15:  neuron_6_mul_27_p <= Pix_771;
    10'd16:  neuron_6_mul_27_p <= Pix_772;
    10'd17:  neuron_6_mul_27_p <= Pix_773;
    10'd18:  neuron_6_mul_27_p <= Pix_774;
    10'd19:  neuron_6_mul_27_p <= Pix_775;
    10'd20:  neuron_6_mul_27_p <= Pix_776;
    10'd21:  neuron_6_mul_27_p <= Pix_777;
    10'd22:  neuron_6_mul_27_p <= Pix_778;
    10'd23:  neuron_6_mul_27_p <= Pix_779;
    10'd24:  neuron_6_mul_27_p <= Pix_780;
    10'd25:  neuron_6_mul_27_p <= Pix_781;
    10'd26:  neuron_6_mul_27_p <= Pix_782;
    10'd27:  neuron_6_mul_27_p <= Pix_783;
    default: neuron_6_mul_27_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_0_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_0_p <= Pix_0;
    10'd1:  neuron_7_mul_0_p <= Pix_1;
    10'd2:  neuron_7_mul_0_p <= Pix_2;
    10'd3:  neuron_7_mul_0_p <= Pix_3;
    10'd4:  neuron_7_mul_0_p <= Pix_4;
    10'd5:  neuron_7_mul_0_p <= Pix_5;
    10'd6:  neuron_7_mul_0_p <= Pix_6;
    10'd7:  neuron_7_mul_0_p <= Pix_7;
    10'd8:  neuron_7_mul_0_p <= Pix_8;
    10'd9:  neuron_7_mul_0_p <= Pix_9;
    10'd10:  neuron_7_mul_0_p <= Pix_10;
    10'd11:  neuron_7_mul_0_p <= Pix_11;
    10'd12:  neuron_7_mul_0_p <= Pix_12;
    10'd13:  neuron_7_mul_0_p <= Pix_13;
    10'd14:  neuron_7_mul_0_p <= Pix_14;
    10'd15:  neuron_7_mul_0_p <= Pix_15;
    10'd16:  neuron_7_mul_0_p <= Pix_16;
    10'd17:  neuron_7_mul_0_p <= Pix_17;
    10'd18:  neuron_7_mul_0_p <= Pix_18;
    10'd19:  neuron_7_mul_0_p <= Pix_19;
    10'd20:  neuron_7_mul_0_p <= Pix_20;
    10'd21:  neuron_7_mul_0_p <= Pix_21;
    10'd22:  neuron_7_mul_0_p <= Pix_22;
    10'd23:  neuron_7_mul_0_p <= Pix_23;
    10'd24:  neuron_7_mul_0_p <= Pix_24;
    10'd25:  neuron_7_mul_0_p <= Pix_25;
    10'd26:  neuron_7_mul_0_p <= Pix_26;
    10'd27:  neuron_7_mul_0_p <= Pix_27;
    default: neuron_7_mul_0_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_1_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_1_p <= Pix_28;
    10'd1:  neuron_7_mul_1_p <= Pix_29;
    10'd2:  neuron_7_mul_1_p <= Pix_30;
    10'd3:  neuron_7_mul_1_p <= Pix_31;
    10'd4:  neuron_7_mul_1_p <= Pix_32;
    10'd5:  neuron_7_mul_1_p <= Pix_33;
    10'd6:  neuron_7_mul_1_p <= Pix_34;
    10'd7:  neuron_7_mul_1_p <= Pix_35;
    10'd8:  neuron_7_mul_1_p <= Pix_36;
    10'd9:  neuron_7_mul_1_p <= Pix_37;
    10'd10:  neuron_7_mul_1_p <= Pix_38;
    10'd11:  neuron_7_mul_1_p <= Pix_39;
    10'd12:  neuron_7_mul_1_p <= Pix_40;
    10'd13:  neuron_7_mul_1_p <= Pix_41;
    10'd14:  neuron_7_mul_1_p <= Pix_42;
    10'd15:  neuron_7_mul_1_p <= Pix_43;
    10'd16:  neuron_7_mul_1_p <= Pix_44;
    10'd17:  neuron_7_mul_1_p <= Pix_45;
    10'd18:  neuron_7_mul_1_p <= Pix_46;
    10'd19:  neuron_7_mul_1_p <= Pix_47;
    10'd20:  neuron_7_mul_1_p <= Pix_48;
    10'd21:  neuron_7_mul_1_p <= Pix_49;
    10'd22:  neuron_7_mul_1_p <= Pix_50;
    10'd23:  neuron_7_mul_1_p <= Pix_51;
    10'd24:  neuron_7_mul_1_p <= Pix_52;
    10'd25:  neuron_7_mul_1_p <= Pix_53;
    10'd26:  neuron_7_mul_1_p <= Pix_54;
    10'd27:  neuron_7_mul_1_p <= Pix_55;
    default: neuron_7_mul_1_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_2_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_2_p <= Pix_56;
    10'd1:  neuron_7_mul_2_p <= Pix_57;
    10'd2:  neuron_7_mul_2_p <= Pix_58;
    10'd3:  neuron_7_mul_2_p <= Pix_59;
    10'd4:  neuron_7_mul_2_p <= Pix_60;
    10'd5:  neuron_7_mul_2_p <= Pix_61;
    10'd6:  neuron_7_mul_2_p <= Pix_62;
    10'd7:  neuron_7_mul_2_p <= Pix_63;
    10'd8:  neuron_7_mul_2_p <= Pix_64;
    10'd9:  neuron_7_mul_2_p <= Pix_65;
    10'd10:  neuron_7_mul_2_p <= Pix_66;
    10'd11:  neuron_7_mul_2_p <= Pix_67;
    10'd12:  neuron_7_mul_2_p <= Pix_68;
    10'd13:  neuron_7_mul_2_p <= Pix_69;
    10'd14:  neuron_7_mul_2_p <= Pix_70;
    10'd15:  neuron_7_mul_2_p <= Pix_71;
    10'd16:  neuron_7_mul_2_p <= Pix_72;
    10'd17:  neuron_7_mul_2_p <= Pix_73;
    10'd18:  neuron_7_mul_2_p <= Pix_74;
    10'd19:  neuron_7_mul_2_p <= Pix_75;
    10'd20:  neuron_7_mul_2_p <= Pix_76;
    10'd21:  neuron_7_mul_2_p <= Pix_77;
    10'd22:  neuron_7_mul_2_p <= Pix_78;
    10'd23:  neuron_7_mul_2_p <= Pix_79;
    10'd24:  neuron_7_mul_2_p <= Pix_80;
    10'd25:  neuron_7_mul_2_p <= Pix_81;
    10'd26:  neuron_7_mul_2_p <= Pix_82;
    10'd27:  neuron_7_mul_2_p <= Pix_83;
    default: neuron_7_mul_2_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_3_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_3_p <= Pix_84;
    10'd1:  neuron_7_mul_3_p <= Pix_85;
    10'd2:  neuron_7_mul_3_p <= Pix_86;
    10'd3:  neuron_7_mul_3_p <= Pix_87;
    10'd4:  neuron_7_mul_3_p <= Pix_88;
    10'd5:  neuron_7_mul_3_p <= Pix_89;
    10'd6:  neuron_7_mul_3_p <= Pix_90;
    10'd7:  neuron_7_mul_3_p <= Pix_91;
    10'd8:  neuron_7_mul_3_p <= Pix_92;
    10'd9:  neuron_7_mul_3_p <= Pix_93;
    10'd10:  neuron_7_mul_3_p <= Pix_94;
    10'd11:  neuron_7_mul_3_p <= Pix_95;
    10'd12:  neuron_7_mul_3_p <= Pix_96;
    10'd13:  neuron_7_mul_3_p <= Pix_97;
    10'd14:  neuron_7_mul_3_p <= Pix_98;
    10'd15:  neuron_7_mul_3_p <= Pix_99;
    10'd16:  neuron_7_mul_3_p <= Pix_100;
    10'd17:  neuron_7_mul_3_p <= Pix_101;
    10'd18:  neuron_7_mul_3_p <= Pix_102;
    10'd19:  neuron_7_mul_3_p <= Pix_103;
    10'd20:  neuron_7_mul_3_p <= Pix_104;
    10'd21:  neuron_7_mul_3_p <= Pix_105;
    10'd22:  neuron_7_mul_3_p <= Pix_106;
    10'd23:  neuron_7_mul_3_p <= Pix_107;
    10'd24:  neuron_7_mul_3_p <= Pix_108;
    10'd25:  neuron_7_mul_3_p <= Pix_109;
    10'd26:  neuron_7_mul_3_p <= Pix_110;
    10'd27:  neuron_7_mul_3_p <= Pix_111;
    default: neuron_7_mul_3_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_4_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_4_p <= Pix_112;
    10'd1:  neuron_7_mul_4_p <= Pix_113;
    10'd2:  neuron_7_mul_4_p <= Pix_114;
    10'd3:  neuron_7_mul_4_p <= Pix_115;
    10'd4:  neuron_7_mul_4_p <= Pix_116;
    10'd5:  neuron_7_mul_4_p <= Pix_117;
    10'd6:  neuron_7_mul_4_p <= Pix_118;
    10'd7:  neuron_7_mul_4_p <= Pix_119;
    10'd8:  neuron_7_mul_4_p <= Pix_120;
    10'd9:  neuron_7_mul_4_p <= Pix_121;
    10'd10:  neuron_7_mul_4_p <= Pix_122;
    10'd11:  neuron_7_mul_4_p <= Pix_123;
    10'd12:  neuron_7_mul_4_p <= Pix_124;
    10'd13:  neuron_7_mul_4_p <= Pix_125;
    10'd14:  neuron_7_mul_4_p <= Pix_126;
    10'd15:  neuron_7_mul_4_p <= Pix_127;
    10'd16:  neuron_7_mul_4_p <= Pix_128;
    10'd17:  neuron_7_mul_4_p <= Pix_129;
    10'd18:  neuron_7_mul_4_p <= Pix_130;
    10'd19:  neuron_7_mul_4_p <= Pix_131;
    10'd20:  neuron_7_mul_4_p <= Pix_132;
    10'd21:  neuron_7_mul_4_p <= Pix_133;
    10'd22:  neuron_7_mul_4_p <= Pix_134;
    10'd23:  neuron_7_mul_4_p <= Pix_135;
    10'd24:  neuron_7_mul_4_p <= Pix_136;
    10'd25:  neuron_7_mul_4_p <= Pix_137;
    10'd26:  neuron_7_mul_4_p <= Pix_138;
    10'd27:  neuron_7_mul_4_p <= Pix_139;
    default: neuron_7_mul_4_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_5_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_5_p <= Pix_140;
    10'd1:  neuron_7_mul_5_p <= Pix_141;
    10'd2:  neuron_7_mul_5_p <= Pix_142;
    10'd3:  neuron_7_mul_5_p <= Pix_143;
    10'd4:  neuron_7_mul_5_p <= Pix_144;
    10'd5:  neuron_7_mul_5_p <= Pix_145;
    10'd6:  neuron_7_mul_5_p <= Pix_146;
    10'd7:  neuron_7_mul_5_p <= Pix_147;
    10'd8:  neuron_7_mul_5_p <= Pix_148;
    10'd9:  neuron_7_mul_5_p <= Pix_149;
    10'd10:  neuron_7_mul_5_p <= Pix_150;
    10'd11:  neuron_7_mul_5_p <= Pix_151;
    10'd12:  neuron_7_mul_5_p <= Pix_152;
    10'd13:  neuron_7_mul_5_p <= Pix_153;
    10'd14:  neuron_7_mul_5_p <= Pix_154;
    10'd15:  neuron_7_mul_5_p <= Pix_155;
    10'd16:  neuron_7_mul_5_p <= Pix_156;
    10'd17:  neuron_7_mul_5_p <= Pix_157;
    10'd18:  neuron_7_mul_5_p <= Pix_158;
    10'd19:  neuron_7_mul_5_p <= Pix_159;
    10'd20:  neuron_7_mul_5_p <= Pix_160;
    10'd21:  neuron_7_mul_5_p <= Pix_161;
    10'd22:  neuron_7_mul_5_p <= Pix_162;
    10'd23:  neuron_7_mul_5_p <= Pix_163;
    10'd24:  neuron_7_mul_5_p <= Pix_164;
    10'd25:  neuron_7_mul_5_p <= Pix_165;
    10'd26:  neuron_7_mul_5_p <= Pix_166;
    10'd27:  neuron_7_mul_5_p <= Pix_167;
    default: neuron_7_mul_5_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_6_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_6_p <= Pix_168;
    10'd1:  neuron_7_mul_6_p <= Pix_169;
    10'd2:  neuron_7_mul_6_p <= Pix_170;
    10'd3:  neuron_7_mul_6_p <= Pix_171;
    10'd4:  neuron_7_mul_6_p <= Pix_172;
    10'd5:  neuron_7_mul_6_p <= Pix_173;
    10'd6:  neuron_7_mul_6_p <= Pix_174;
    10'd7:  neuron_7_mul_6_p <= Pix_175;
    10'd8:  neuron_7_mul_6_p <= Pix_176;
    10'd9:  neuron_7_mul_6_p <= Pix_177;
    10'd10:  neuron_7_mul_6_p <= Pix_178;
    10'd11:  neuron_7_mul_6_p <= Pix_179;
    10'd12:  neuron_7_mul_6_p <= Pix_180;
    10'd13:  neuron_7_mul_6_p <= Pix_181;
    10'd14:  neuron_7_mul_6_p <= Pix_182;
    10'd15:  neuron_7_mul_6_p <= Pix_183;
    10'd16:  neuron_7_mul_6_p <= Pix_184;
    10'd17:  neuron_7_mul_6_p <= Pix_185;
    10'd18:  neuron_7_mul_6_p <= Pix_186;
    10'd19:  neuron_7_mul_6_p <= Pix_187;
    10'd20:  neuron_7_mul_6_p <= Pix_188;
    10'd21:  neuron_7_mul_6_p <= Pix_189;
    10'd22:  neuron_7_mul_6_p <= Pix_190;
    10'd23:  neuron_7_mul_6_p <= Pix_191;
    10'd24:  neuron_7_mul_6_p <= Pix_192;
    10'd25:  neuron_7_mul_6_p <= Pix_193;
    10'd26:  neuron_7_mul_6_p <= Pix_194;
    10'd27:  neuron_7_mul_6_p <= Pix_195;
    default: neuron_7_mul_6_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_7_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_7_p <= Pix_196;
    10'd1:  neuron_7_mul_7_p <= Pix_197;
    10'd2:  neuron_7_mul_7_p <= Pix_198;
    10'd3:  neuron_7_mul_7_p <= Pix_199;
    10'd4:  neuron_7_mul_7_p <= Pix_200;
    10'd5:  neuron_7_mul_7_p <= Pix_201;
    10'd6:  neuron_7_mul_7_p <= Pix_202;
    10'd7:  neuron_7_mul_7_p <= Pix_203;
    10'd8:  neuron_7_mul_7_p <= Pix_204;
    10'd9:  neuron_7_mul_7_p <= Pix_205;
    10'd10:  neuron_7_mul_7_p <= Pix_206;
    10'd11:  neuron_7_mul_7_p <= Pix_207;
    10'd12:  neuron_7_mul_7_p <= Pix_208;
    10'd13:  neuron_7_mul_7_p <= Pix_209;
    10'd14:  neuron_7_mul_7_p <= Pix_210;
    10'd15:  neuron_7_mul_7_p <= Pix_211;
    10'd16:  neuron_7_mul_7_p <= Pix_212;
    10'd17:  neuron_7_mul_7_p <= Pix_213;
    10'd18:  neuron_7_mul_7_p <= Pix_214;
    10'd19:  neuron_7_mul_7_p <= Pix_215;
    10'd20:  neuron_7_mul_7_p <= Pix_216;
    10'd21:  neuron_7_mul_7_p <= Pix_217;
    10'd22:  neuron_7_mul_7_p <= Pix_218;
    10'd23:  neuron_7_mul_7_p <= Pix_219;
    10'd24:  neuron_7_mul_7_p <= Pix_220;
    10'd25:  neuron_7_mul_7_p <= Pix_221;
    10'd26:  neuron_7_mul_7_p <= Pix_222;
    10'd27:  neuron_7_mul_7_p <= Pix_223;
    default: neuron_7_mul_7_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_8_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_8_p <= Pix_224;
    10'd1:  neuron_7_mul_8_p <= Pix_225;
    10'd2:  neuron_7_mul_8_p <= Pix_226;
    10'd3:  neuron_7_mul_8_p <= Pix_227;
    10'd4:  neuron_7_mul_8_p <= Pix_228;
    10'd5:  neuron_7_mul_8_p <= Pix_229;
    10'd6:  neuron_7_mul_8_p <= Pix_230;
    10'd7:  neuron_7_mul_8_p <= Pix_231;
    10'd8:  neuron_7_mul_8_p <= Pix_232;
    10'd9:  neuron_7_mul_8_p <= Pix_233;
    10'd10:  neuron_7_mul_8_p <= Pix_234;
    10'd11:  neuron_7_mul_8_p <= Pix_235;
    10'd12:  neuron_7_mul_8_p <= Pix_236;
    10'd13:  neuron_7_mul_8_p <= Pix_237;
    10'd14:  neuron_7_mul_8_p <= Pix_238;
    10'd15:  neuron_7_mul_8_p <= Pix_239;
    10'd16:  neuron_7_mul_8_p <= Pix_240;
    10'd17:  neuron_7_mul_8_p <= Pix_241;
    10'd18:  neuron_7_mul_8_p <= Pix_242;
    10'd19:  neuron_7_mul_8_p <= Pix_243;
    10'd20:  neuron_7_mul_8_p <= Pix_244;
    10'd21:  neuron_7_mul_8_p <= Pix_245;
    10'd22:  neuron_7_mul_8_p <= Pix_246;
    10'd23:  neuron_7_mul_8_p <= Pix_247;
    10'd24:  neuron_7_mul_8_p <= Pix_248;
    10'd25:  neuron_7_mul_8_p <= Pix_249;
    10'd26:  neuron_7_mul_8_p <= Pix_250;
    10'd27:  neuron_7_mul_8_p <= Pix_251;
    default: neuron_7_mul_8_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_9_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_9_p <= Pix_252;
    10'd1:  neuron_7_mul_9_p <= Pix_253;
    10'd2:  neuron_7_mul_9_p <= Pix_254;
    10'd3:  neuron_7_mul_9_p <= Pix_255;
    10'd4:  neuron_7_mul_9_p <= Pix_256;
    10'd5:  neuron_7_mul_9_p <= Pix_257;
    10'd6:  neuron_7_mul_9_p <= Pix_258;
    10'd7:  neuron_7_mul_9_p <= Pix_259;
    10'd8:  neuron_7_mul_9_p <= Pix_260;
    10'd9:  neuron_7_mul_9_p <= Pix_261;
    10'd10:  neuron_7_mul_9_p <= Pix_262;
    10'd11:  neuron_7_mul_9_p <= Pix_263;
    10'd12:  neuron_7_mul_9_p <= Pix_264;
    10'd13:  neuron_7_mul_9_p <= Pix_265;
    10'd14:  neuron_7_mul_9_p <= Pix_266;
    10'd15:  neuron_7_mul_9_p <= Pix_267;
    10'd16:  neuron_7_mul_9_p <= Pix_268;
    10'd17:  neuron_7_mul_9_p <= Pix_269;
    10'd18:  neuron_7_mul_9_p <= Pix_270;
    10'd19:  neuron_7_mul_9_p <= Pix_271;
    10'd20:  neuron_7_mul_9_p <= Pix_272;
    10'd21:  neuron_7_mul_9_p <= Pix_273;
    10'd22:  neuron_7_mul_9_p <= Pix_274;
    10'd23:  neuron_7_mul_9_p <= Pix_275;
    10'd24:  neuron_7_mul_9_p <= Pix_276;
    10'd25:  neuron_7_mul_9_p <= Pix_277;
    10'd26:  neuron_7_mul_9_p <= Pix_278;
    10'd27:  neuron_7_mul_9_p <= Pix_279;
    default: neuron_7_mul_9_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_10_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_10_p <= Pix_280;
    10'd1:  neuron_7_mul_10_p <= Pix_281;
    10'd2:  neuron_7_mul_10_p <= Pix_282;
    10'd3:  neuron_7_mul_10_p <= Pix_283;
    10'd4:  neuron_7_mul_10_p <= Pix_284;
    10'd5:  neuron_7_mul_10_p <= Pix_285;
    10'd6:  neuron_7_mul_10_p <= Pix_286;
    10'd7:  neuron_7_mul_10_p <= Pix_287;
    10'd8:  neuron_7_mul_10_p <= Pix_288;
    10'd9:  neuron_7_mul_10_p <= Pix_289;
    10'd10:  neuron_7_mul_10_p <= Pix_290;
    10'd11:  neuron_7_mul_10_p <= Pix_291;
    10'd12:  neuron_7_mul_10_p <= Pix_292;
    10'd13:  neuron_7_mul_10_p <= Pix_293;
    10'd14:  neuron_7_mul_10_p <= Pix_294;
    10'd15:  neuron_7_mul_10_p <= Pix_295;
    10'd16:  neuron_7_mul_10_p <= Pix_296;
    10'd17:  neuron_7_mul_10_p <= Pix_297;
    10'd18:  neuron_7_mul_10_p <= Pix_298;
    10'd19:  neuron_7_mul_10_p <= Pix_299;
    10'd20:  neuron_7_mul_10_p <= Pix_300;
    10'd21:  neuron_7_mul_10_p <= Pix_301;
    10'd22:  neuron_7_mul_10_p <= Pix_302;
    10'd23:  neuron_7_mul_10_p <= Pix_303;
    10'd24:  neuron_7_mul_10_p <= Pix_304;
    10'd25:  neuron_7_mul_10_p <= Pix_305;
    10'd26:  neuron_7_mul_10_p <= Pix_306;
    10'd27:  neuron_7_mul_10_p <= Pix_307;
    default: neuron_7_mul_10_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_11_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_11_p <= Pix_308;
    10'd1:  neuron_7_mul_11_p <= Pix_309;
    10'd2:  neuron_7_mul_11_p <= Pix_310;
    10'd3:  neuron_7_mul_11_p <= Pix_311;
    10'd4:  neuron_7_mul_11_p <= Pix_312;
    10'd5:  neuron_7_mul_11_p <= Pix_313;
    10'd6:  neuron_7_mul_11_p <= Pix_314;
    10'd7:  neuron_7_mul_11_p <= Pix_315;
    10'd8:  neuron_7_mul_11_p <= Pix_316;
    10'd9:  neuron_7_mul_11_p <= Pix_317;
    10'd10:  neuron_7_mul_11_p <= Pix_318;
    10'd11:  neuron_7_mul_11_p <= Pix_319;
    10'd12:  neuron_7_mul_11_p <= Pix_320;
    10'd13:  neuron_7_mul_11_p <= Pix_321;
    10'd14:  neuron_7_mul_11_p <= Pix_322;
    10'd15:  neuron_7_mul_11_p <= Pix_323;
    10'd16:  neuron_7_mul_11_p <= Pix_324;
    10'd17:  neuron_7_mul_11_p <= Pix_325;
    10'd18:  neuron_7_mul_11_p <= Pix_326;
    10'd19:  neuron_7_mul_11_p <= Pix_327;
    10'd20:  neuron_7_mul_11_p <= Pix_328;
    10'd21:  neuron_7_mul_11_p <= Pix_329;
    10'd22:  neuron_7_mul_11_p <= Pix_330;
    10'd23:  neuron_7_mul_11_p <= Pix_331;
    10'd24:  neuron_7_mul_11_p <= Pix_332;
    10'd25:  neuron_7_mul_11_p <= Pix_333;
    10'd26:  neuron_7_mul_11_p <= Pix_334;
    10'd27:  neuron_7_mul_11_p <= Pix_335;
    default: neuron_7_mul_11_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_12_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_12_p <= Pix_336;
    10'd1:  neuron_7_mul_12_p <= Pix_337;
    10'd2:  neuron_7_mul_12_p <= Pix_338;
    10'd3:  neuron_7_mul_12_p <= Pix_339;
    10'd4:  neuron_7_mul_12_p <= Pix_340;
    10'd5:  neuron_7_mul_12_p <= Pix_341;
    10'd6:  neuron_7_mul_12_p <= Pix_342;
    10'd7:  neuron_7_mul_12_p <= Pix_343;
    10'd8:  neuron_7_mul_12_p <= Pix_344;
    10'd9:  neuron_7_mul_12_p <= Pix_345;
    10'd10:  neuron_7_mul_12_p <= Pix_346;
    10'd11:  neuron_7_mul_12_p <= Pix_347;
    10'd12:  neuron_7_mul_12_p <= Pix_348;
    10'd13:  neuron_7_mul_12_p <= Pix_349;
    10'd14:  neuron_7_mul_12_p <= Pix_350;
    10'd15:  neuron_7_mul_12_p <= Pix_351;
    10'd16:  neuron_7_mul_12_p <= Pix_352;
    10'd17:  neuron_7_mul_12_p <= Pix_353;
    10'd18:  neuron_7_mul_12_p <= Pix_354;
    10'd19:  neuron_7_mul_12_p <= Pix_355;
    10'd20:  neuron_7_mul_12_p <= Pix_356;
    10'd21:  neuron_7_mul_12_p <= Pix_357;
    10'd22:  neuron_7_mul_12_p <= Pix_358;
    10'd23:  neuron_7_mul_12_p <= Pix_359;
    10'd24:  neuron_7_mul_12_p <= Pix_360;
    10'd25:  neuron_7_mul_12_p <= Pix_361;
    10'd26:  neuron_7_mul_12_p <= Pix_362;
    10'd27:  neuron_7_mul_12_p <= Pix_363;
    default: neuron_7_mul_12_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_13_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_13_p <= Pix_364;
    10'd1:  neuron_7_mul_13_p <= Pix_365;
    10'd2:  neuron_7_mul_13_p <= Pix_366;
    10'd3:  neuron_7_mul_13_p <= Pix_367;
    10'd4:  neuron_7_mul_13_p <= Pix_368;
    10'd5:  neuron_7_mul_13_p <= Pix_369;
    10'd6:  neuron_7_mul_13_p <= Pix_370;
    10'd7:  neuron_7_mul_13_p <= Pix_371;
    10'd8:  neuron_7_mul_13_p <= Pix_372;
    10'd9:  neuron_7_mul_13_p <= Pix_373;
    10'd10:  neuron_7_mul_13_p <= Pix_374;
    10'd11:  neuron_7_mul_13_p <= Pix_375;
    10'd12:  neuron_7_mul_13_p <= Pix_376;
    10'd13:  neuron_7_mul_13_p <= Pix_377;
    10'd14:  neuron_7_mul_13_p <= Pix_378;
    10'd15:  neuron_7_mul_13_p <= Pix_379;
    10'd16:  neuron_7_mul_13_p <= Pix_380;
    10'd17:  neuron_7_mul_13_p <= Pix_381;
    10'd18:  neuron_7_mul_13_p <= Pix_382;
    10'd19:  neuron_7_mul_13_p <= Pix_383;
    10'd20:  neuron_7_mul_13_p <= Pix_384;
    10'd21:  neuron_7_mul_13_p <= Pix_385;
    10'd22:  neuron_7_mul_13_p <= Pix_386;
    10'd23:  neuron_7_mul_13_p <= Pix_387;
    10'd24:  neuron_7_mul_13_p <= Pix_388;
    10'd25:  neuron_7_mul_13_p <= Pix_389;
    10'd26:  neuron_7_mul_13_p <= Pix_390;
    10'd27:  neuron_7_mul_13_p <= Pix_391;
    default: neuron_7_mul_13_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_14_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_14_p <= Pix_392;
    10'd1:  neuron_7_mul_14_p <= Pix_393;
    10'd2:  neuron_7_mul_14_p <= Pix_394;
    10'd3:  neuron_7_mul_14_p <= Pix_395;
    10'd4:  neuron_7_mul_14_p <= Pix_396;
    10'd5:  neuron_7_mul_14_p <= Pix_397;
    10'd6:  neuron_7_mul_14_p <= Pix_398;
    10'd7:  neuron_7_mul_14_p <= Pix_399;
    10'd8:  neuron_7_mul_14_p <= Pix_400;
    10'd9:  neuron_7_mul_14_p <= Pix_401;
    10'd10:  neuron_7_mul_14_p <= Pix_402;
    10'd11:  neuron_7_mul_14_p <= Pix_403;
    10'd12:  neuron_7_mul_14_p <= Pix_404;
    10'd13:  neuron_7_mul_14_p <= Pix_405;
    10'd14:  neuron_7_mul_14_p <= Pix_406;
    10'd15:  neuron_7_mul_14_p <= Pix_407;
    10'd16:  neuron_7_mul_14_p <= Pix_408;
    10'd17:  neuron_7_mul_14_p <= Pix_409;
    10'd18:  neuron_7_mul_14_p <= Pix_410;
    10'd19:  neuron_7_mul_14_p <= Pix_411;
    10'd20:  neuron_7_mul_14_p <= Pix_412;
    10'd21:  neuron_7_mul_14_p <= Pix_413;
    10'd22:  neuron_7_mul_14_p <= Pix_414;
    10'd23:  neuron_7_mul_14_p <= Pix_415;
    10'd24:  neuron_7_mul_14_p <= Pix_416;
    10'd25:  neuron_7_mul_14_p <= Pix_417;
    10'd26:  neuron_7_mul_14_p <= Pix_418;
    10'd27:  neuron_7_mul_14_p <= Pix_419;
    default: neuron_7_mul_14_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_15_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_15_p <= Pix_420;
    10'd1:  neuron_7_mul_15_p <= Pix_421;
    10'd2:  neuron_7_mul_15_p <= Pix_422;
    10'd3:  neuron_7_mul_15_p <= Pix_423;
    10'd4:  neuron_7_mul_15_p <= Pix_424;
    10'd5:  neuron_7_mul_15_p <= Pix_425;
    10'd6:  neuron_7_mul_15_p <= Pix_426;
    10'd7:  neuron_7_mul_15_p <= Pix_427;
    10'd8:  neuron_7_mul_15_p <= Pix_428;
    10'd9:  neuron_7_mul_15_p <= Pix_429;
    10'd10:  neuron_7_mul_15_p <= Pix_430;
    10'd11:  neuron_7_mul_15_p <= Pix_431;
    10'd12:  neuron_7_mul_15_p <= Pix_432;
    10'd13:  neuron_7_mul_15_p <= Pix_433;
    10'd14:  neuron_7_mul_15_p <= Pix_434;
    10'd15:  neuron_7_mul_15_p <= Pix_435;
    10'd16:  neuron_7_mul_15_p <= Pix_436;
    10'd17:  neuron_7_mul_15_p <= Pix_437;
    10'd18:  neuron_7_mul_15_p <= Pix_438;
    10'd19:  neuron_7_mul_15_p <= Pix_439;
    10'd20:  neuron_7_mul_15_p <= Pix_440;
    10'd21:  neuron_7_mul_15_p <= Pix_441;
    10'd22:  neuron_7_mul_15_p <= Pix_442;
    10'd23:  neuron_7_mul_15_p <= Pix_443;
    10'd24:  neuron_7_mul_15_p <= Pix_444;
    10'd25:  neuron_7_mul_15_p <= Pix_445;
    10'd26:  neuron_7_mul_15_p <= Pix_446;
    10'd27:  neuron_7_mul_15_p <= Pix_447;
    default: neuron_7_mul_15_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_16_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_16_p <= Pix_448;
    10'd1:  neuron_7_mul_16_p <= Pix_449;
    10'd2:  neuron_7_mul_16_p <= Pix_450;
    10'd3:  neuron_7_mul_16_p <= Pix_451;
    10'd4:  neuron_7_mul_16_p <= Pix_452;
    10'd5:  neuron_7_mul_16_p <= Pix_453;
    10'd6:  neuron_7_mul_16_p <= Pix_454;
    10'd7:  neuron_7_mul_16_p <= Pix_455;
    10'd8:  neuron_7_mul_16_p <= Pix_456;
    10'd9:  neuron_7_mul_16_p <= Pix_457;
    10'd10:  neuron_7_mul_16_p <= Pix_458;
    10'd11:  neuron_7_mul_16_p <= Pix_459;
    10'd12:  neuron_7_mul_16_p <= Pix_460;
    10'd13:  neuron_7_mul_16_p <= Pix_461;
    10'd14:  neuron_7_mul_16_p <= Pix_462;
    10'd15:  neuron_7_mul_16_p <= Pix_463;
    10'd16:  neuron_7_mul_16_p <= Pix_464;
    10'd17:  neuron_7_mul_16_p <= Pix_465;
    10'd18:  neuron_7_mul_16_p <= Pix_466;
    10'd19:  neuron_7_mul_16_p <= Pix_467;
    10'd20:  neuron_7_mul_16_p <= Pix_468;
    10'd21:  neuron_7_mul_16_p <= Pix_469;
    10'd22:  neuron_7_mul_16_p <= Pix_470;
    10'd23:  neuron_7_mul_16_p <= Pix_471;
    10'd24:  neuron_7_mul_16_p <= Pix_472;
    10'd25:  neuron_7_mul_16_p <= Pix_473;
    10'd26:  neuron_7_mul_16_p <= Pix_474;
    10'd27:  neuron_7_mul_16_p <= Pix_475;
    default: neuron_7_mul_16_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_17_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_17_p <= Pix_476;
    10'd1:  neuron_7_mul_17_p <= Pix_477;
    10'd2:  neuron_7_mul_17_p <= Pix_478;
    10'd3:  neuron_7_mul_17_p <= Pix_479;
    10'd4:  neuron_7_mul_17_p <= Pix_480;
    10'd5:  neuron_7_mul_17_p <= Pix_481;
    10'd6:  neuron_7_mul_17_p <= Pix_482;
    10'd7:  neuron_7_mul_17_p <= Pix_483;
    10'd8:  neuron_7_mul_17_p <= Pix_484;
    10'd9:  neuron_7_mul_17_p <= Pix_485;
    10'd10:  neuron_7_mul_17_p <= Pix_486;
    10'd11:  neuron_7_mul_17_p <= Pix_487;
    10'd12:  neuron_7_mul_17_p <= Pix_488;
    10'd13:  neuron_7_mul_17_p <= Pix_489;
    10'd14:  neuron_7_mul_17_p <= Pix_490;
    10'd15:  neuron_7_mul_17_p <= Pix_491;
    10'd16:  neuron_7_mul_17_p <= Pix_492;
    10'd17:  neuron_7_mul_17_p <= Pix_493;
    10'd18:  neuron_7_mul_17_p <= Pix_494;
    10'd19:  neuron_7_mul_17_p <= Pix_495;
    10'd20:  neuron_7_mul_17_p <= Pix_496;
    10'd21:  neuron_7_mul_17_p <= Pix_497;
    10'd22:  neuron_7_mul_17_p <= Pix_498;
    10'd23:  neuron_7_mul_17_p <= Pix_499;
    10'd24:  neuron_7_mul_17_p <= Pix_500;
    10'd25:  neuron_7_mul_17_p <= Pix_501;
    10'd26:  neuron_7_mul_17_p <= Pix_502;
    10'd27:  neuron_7_mul_17_p <= Pix_503;
    default: neuron_7_mul_17_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_18_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_18_p <= Pix_504;
    10'd1:  neuron_7_mul_18_p <= Pix_505;
    10'd2:  neuron_7_mul_18_p <= Pix_506;
    10'd3:  neuron_7_mul_18_p <= Pix_507;
    10'd4:  neuron_7_mul_18_p <= Pix_508;
    10'd5:  neuron_7_mul_18_p <= Pix_509;
    10'd6:  neuron_7_mul_18_p <= Pix_510;
    10'd7:  neuron_7_mul_18_p <= Pix_511;
    10'd8:  neuron_7_mul_18_p <= Pix_512;
    10'd9:  neuron_7_mul_18_p <= Pix_513;
    10'd10:  neuron_7_mul_18_p <= Pix_514;
    10'd11:  neuron_7_mul_18_p <= Pix_515;
    10'd12:  neuron_7_mul_18_p <= Pix_516;
    10'd13:  neuron_7_mul_18_p <= Pix_517;
    10'd14:  neuron_7_mul_18_p <= Pix_518;
    10'd15:  neuron_7_mul_18_p <= Pix_519;
    10'd16:  neuron_7_mul_18_p <= Pix_520;
    10'd17:  neuron_7_mul_18_p <= Pix_521;
    10'd18:  neuron_7_mul_18_p <= Pix_522;
    10'd19:  neuron_7_mul_18_p <= Pix_523;
    10'd20:  neuron_7_mul_18_p <= Pix_524;
    10'd21:  neuron_7_mul_18_p <= Pix_525;
    10'd22:  neuron_7_mul_18_p <= Pix_526;
    10'd23:  neuron_7_mul_18_p <= Pix_527;
    10'd24:  neuron_7_mul_18_p <= Pix_528;
    10'd25:  neuron_7_mul_18_p <= Pix_529;
    10'd26:  neuron_7_mul_18_p <= Pix_530;
    10'd27:  neuron_7_mul_18_p <= Pix_531;
    default: neuron_7_mul_18_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_19_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_19_p <= Pix_532;
    10'd1:  neuron_7_mul_19_p <= Pix_533;
    10'd2:  neuron_7_mul_19_p <= Pix_534;
    10'd3:  neuron_7_mul_19_p <= Pix_535;
    10'd4:  neuron_7_mul_19_p <= Pix_536;
    10'd5:  neuron_7_mul_19_p <= Pix_537;
    10'd6:  neuron_7_mul_19_p <= Pix_538;
    10'd7:  neuron_7_mul_19_p <= Pix_539;
    10'd8:  neuron_7_mul_19_p <= Pix_540;
    10'd9:  neuron_7_mul_19_p <= Pix_541;
    10'd10:  neuron_7_mul_19_p <= Pix_542;
    10'd11:  neuron_7_mul_19_p <= Pix_543;
    10'd12:  neuron_7_mul_19_p <= Pix_544;
    10'd13:  neuron_7_mul_19_p <= Pix_545;
    10'd14:  neuron_7_mul_19_p <= Pix_546;
    10'd15:  neuron_7_mul_19_p <= Pix_547;
    10'd16:  neuron_7_mul_19_p <= Pix_548;
    10'd17:  neuron_7_mul_19_p <= Pix_549;
    10'd18:  neuron_7_mul_19_p <= Pix_550;
    10'd19:  neuron_7_mul_19_p <= Pix_551;
    10'd20:  neuron_7_mul_19_p <= Pix_552;
    10'd21:  neuron_7_mul_19_p <= Pix_553;
    10'd22:  neuron_7_mul_19_p <= Pix_554;
    10'd23:  neuron_7_mul_19_p <= Pix_555;
    10'd24:  neuron_7_mul_19_p <= Pix_556;
    10'd25:  neuron_7_mul_19_p <= Pix_557;
    10'd26:  neuron_7_mul_19_p <= Pix_558;
    10'd27:  neuron_7_mul_19_p <= Pix_559;
    default: neuron_7_mul_19_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_20_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_20_p <= Pix_560;
    10'd1:  neuron_7_mul_20_p <= Pix_561;
    10'd2:  neuron_7_mul_20_p <= Pix_562;
    10'd3:  neuron_7_mul_20_p <= Pix_563;
    10'd4:  neuron_7_mul_20_p <= Pix_564;
    10'd5:  neuron_7_mul_20_p <= Pix_565;
    10'd6:  neuron_7_mul_20_p <= Pix_566;
    10'd7:  neuron_7_mul_20_p <= Pix_567;
    10'd8:  neuron_7_mul_20_p <= Pix_568;
    10'd9:  neuron_7_mul_20_p <= Pix_569;
    10'd10:  neuron_7_mul_20_p <= Pix_570;
    10'd11:  neuron_7_mul_20_p <= Pix_571;
    10'd12:  neuron_7_mul_20_p <= Pix_572;
    10'd13:  neuron_7_mul_20_p <= Pix_573;
    10'd14:  neuron_7_mul_20_p <= Pix_574;
    10'd15:  neuron_7_mul_20_p <= Pix_575;
    10'd16:  neuron_7_mul_20_p <= Pix_576;
    10'd17:  neuron_7_mul_20_p <= Pix_577;
    10'd18:  neuron_7_mul_20_p <= Pix_578;
    10'd19:  neuron_7_mul_20_p <= Pix_579;
    10'd20:  neuron_7_mul_20_p <= Pix_580;
    10'd21:  neuron_7_mul_20_p <= Pix_581;
    10'd22:  neuron_7_mul_20_p <= Pix_582;
    10'd23:  neuron_7_mul_20_p <= Pix_583;
    10'd24:  neuron_7_mul_20_p <= Pix_584;
    10'd25:  neuron_7_mul_20_p <= Pix_585;
    10'd26:  neuron_7_mul_20_p <= Pix_586;
    10'd27:  neuron_7_mul_20_p <= Pix_587;
    default: neuron_7_mul_20_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_21_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_21_p <= Pix_588;
    10'd1:  neuron_7_mul_21_p <= Pix_589;
    10'd2:  neuron_7_mul_21_p <= Pix_590;
    10'd3:  neuron_7_mul_21_p <= Pix_591;
    10'd4:  neuron_7_mul_21_p <= Pix_592;
    10'd5:  neuron_7_mul_21_p <= Pix_593;
    10'd6:  neuron_7_mul_21_p <= Pix_594;
    10'd7:  neuron_7_mul_21_p <= Pix_595;
    10'd8:  neuron_7_mul_21_p <= Pix_596;
    10'd9:  neuron_7_mul_21_p <= Pix_597;
    10'd10:  neuron_7_mul_21_p <= Pix_598;
    10'd11:  neuron_7_mul_21_p <= Pix_599;
    10'd12:  neuron_7_mul_21_p <= Pix_600;
    10'd13:  neuron_7_mul_21_p <= Pix_601;
    10'd14:  neuron_7_mul_21_p <= Pix_602;
    10'd15:  neuron_7_mul_21_p <= Pix_603;
    10'd16:  neuron_7_mul_21_p <= Pix_604;
    10'd17:  neuron_7_mul_21_p <= Pix_605;
    10'd18:  neuron_7_mul_21_p <= Pix_606;
    10'd19:  neuron_7_mul_21_p <= Pix_607;
    10'd20:  neuron_7_mul_21_p <= Pix_608;
    10'd21:  neuron_7_mul_21_p <= Pix_609;
    10'd22:  neuron_7_mul_21_p <= Pix_610;
    10'd23:  neuron_7_mul_21_p <= Pix_611;
    10'd24:  neuron_7_mul_21_p <= Pix_612;
    10'd25:  neuron_7_mul_21_p <= Pix_613;
    10'd26:  neuron_7_mul_21_p <= Pix_614;
    10'd27:  neuron_7_mul_21_p <= Pix_615;
    default: neuron_7_mul_21_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_22_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_22_p <= Pix_616;
    10'd1:  neuron_7_mul_22_p <= Pix_617;
    10'd2:  neuron_7_mul_22_p <= Pix_618;
    10'd3:  neuron_7_mul_22_p <= Pix_619;
    10'd4:  neuron_7_mul_22_p <= Pix_620;
    10'd5:  neuron_7_mul_22_p <= Pix_621;
    10'd6:  neuron_7_mul_22_p <= Pix_622;
    10'd7:  neuron_7_mul_22_p <= Pix_623;
    10'd8:  neuron_7_mul_22_p <= Pix_624;
    10'd9:  neuron_7_mul_22_p <= Pix_625;
    10'd10:  neuron_7_mul_22_p <= Pix_626;
    10'd11:  neuron_7_mul_22_p <= Pix_627;
    10'd12:  neuron_7_mul_22_p <= Pix_628;
    10'd13:  neuron_7_mul_22_p <= Pix_629;
    10'd14:  neuron_7_mul_22_p <= Pix_630;
    10'd15:  neuron_7_mul_22_p <= Pix_631;
    10'd16:  neuron_7_mul_22_p <= Pix_632;
    10'd17:  neuron_7_mul_22_p <= Pix_633;
    10'd18:  neuron_7_mul_22_p <= Pix_634;
    10'd19:  neuron_7_mul_22_p <= Pix_635;
    10'd20:  neuron_7_mul_22_p <= Pix_636;
    10'd21:  neuron_7_mul_22_p <= Pix_637;
    10'd22:  neuron_7_mul_22_p <= Pix_638;
    10'd23:  neuron_7_mul_22_p <= Pix_639;
    10'd24:  neuron_7_mul_22_p <= Pix_640;
    10'd25:  neuron_7_mul_22_p <= Pix_641;
    10'd26:  neuron_7_mul_22_p <= Pix_642;
    10'd27:  neuron_7_mul_22_p <= Pix_643;
    default: neuron_7_mul_22_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_23_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_23_p <= Pix_644;
    10'd1:  neuron_7_mul_23_p <= Pix_645;
    10'd2:  neuron_7_mul_23_p <= Pix_646;
    10'd3:  neuron_7_mul_23_p <= Pix_647;
    10'd4:  neuron_7_mul_23_p <= Pix_648;
    10'd5:  neuron_7_mul_23_p <= Pix_649;
    10'd6:  neuron_7_mul_23_p <= Pix_650;
    10'd7:  neuron_7_mul_23_p <= Pix_651;
    10'd8:  neuron_7_mul_23_p <= Pix_652;
    10'd9:  neuron_7_mul_23_p <= Pix_653;
    10'd10:  neuron_7_mul_23_p <= Pix_654;
    10'd11:  neuron_7_mul_23_p <= Pix_655;
    10'd12:  neuron_7_mul_23_p <= Pix_656;
    10'd13:  neuron_7_mul_23_p <= Pix_657;
    10'd14:  neuron_7_mul_23_p <= Pix_658;
    10'd15:  neuron_7_mul_23_p <= Pix_659;
    10'd16:  neuron_7_mul_23_p <= Pix_660;
    10'd17:  neuron_7_mul_23_p <= Pix_661;
    10'd18:  neuron_7_mul_23_p <= Pix_662;
    10'd19:  neuron_7_mul_23_p <= Pix_663;
    10'd20:  neuron_7_mul_23_p <= Pix_664;
    10'd21:  neuron_7_mul_23_p <= Pix_665;
    10'd22:  neuron_7_mul_23_p <= Pix_666;
    10'd23:  neuron_7_mul_23_p <= Pix_667;
    10'd24:  neuron_7_mul_23_p <= Pix_668;
    10'd25:  neuron_7_mul_23_p <= Pix_669;
    10'd26:  neuron_7_mul_23_p <= Pix_670;
    10'd27:  neuron_7_mul_23_p <= Pix_671;
    default: neuron_7_mul_23_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_24_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_24_p <= Pix_672;
    10'd1:  neuron_7_mul_24_p <= Pix_673;
    10'd2:  neuron_7_mul_24_p <= Pix_674;
    10'd3:  neuron_7_mul_24_p <= Pix_675;
    10'd4:  neuron_7_mul_24_p <= Pix_676;
    10'd5:  neuron_7_mul_24_p <= Pix_677;
    10'd6:  neuron_7_mul_24_p <= Pix_678;
    10'd7:  neuron_7_mul_24_p <= Pix_679;
    10'd8:  neuron_7_mul_24_p <= Pix_680;
    10'd9:  neuron_7_mul_24_p <= Pix_681;
    10'd10:  neuron_7_mul_24_p <= Pix_682;
    10'd11:  neuron_7_mul_24_p <= Pix_683;
    10'd12:  neuron_7_mul_24_p <= Pix_684;
    10'd13:  neuron_7_mul_24_p <= Pix_685;
    10'd14:  neuron_7_mul_24_p <= Pix_686;
    10'd15:  neuron_7_mul_24_p <= Pix_687;
    10'd16:  neuron_7_mul_24_p <= Pix_688;
    10'd17:  neuron_7_mul_24_p <= Pix_689;
    10'd18:  neuron_7_mul_24_p <= Pix_690;
    10'd19:  neuron_7_mul_24_p <= Pix_691;
    10'd20:  neuron_7_mul_24_p <= Pix_692;
    10'd21:  neuron_7_mul_24_p <= Pix_693;
    10'd22:  neuron_7_mul_24_p <= Pix_694;
    10'd23:  neuron_7_mul_24_p <= Pix_695;
    10'd24:  neuron_7_mul_24_p <= Pix_696;
    10'd25:  neuron_7_mul_24_p <= Pix_697;
    10'd26:  neuron_7_mul_24_p <= Pix_698;
    10'd27:  neuron_7_mul_24_p <= Pix_699;
    default: neuron_7_mul_24_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_25_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_25_p <= Pix_700;
    10'd1:  neuron_7_mul_25_p <= Pix_701;
    10'd2:  neuron_7_mul_25_p <= Pix_702;
    10'd3:  neuron_7_mul_25_p <= Pix_703;
    10'd4:  neuron_7_mul_25_p <= Pix_704;
    10'd5:  neuron_7_mul_25_p <= Pix_705;
    10'd6:  neuron_7_mul_25_p <= Pix_706;
    10'd7:  neuron_7_mul_25_p <= Pix_707;
    10'd8:  neuron_7_mul_25_p <= Pix_708;
    10'd9:  neuron_7_mul_25_p <= Pix_709;
    10'd10:  neuron_7_mul_25_p <= Pix_710;
    10'd11:  neuron_7_mul_25_p <= Pix_711;
    10'd12:  neuron_7_mul_25_p <= Pix_712;
    10'd13:  neuron_7_mul_25_p <= Pix_713;
    10'd14:  neuron_7_mul_25_p <= Pix_714;
    10'd15:  neuron_7_mul_25_p <= Pix_715;
    10'd16:  neuron_7_mul_25_p <= Pix_716;
    10'd17:  neuron_7_mul_25_p <= Pix_717;
    10'd18:  neuron_7_mul_25_p <= Pix_718;
    10'd19:  neuron_7_mul_25_p <= Pix_719;
    10'd20:  neuron_7_mul_25_p <= Pix_720;
    10'd21:  neuron_7_mul_25_p <= Pix_721;
    10'd22:  neuron_7_mul_25_p <= Pix_722;
    10'd23:  neuron_7_mul_25_p <= Pix_723;
    10'd24:  neuron_7_mul_25_p <= Pix_724;
    10'd25:  neuron_7_mul_25_p <= Pix_725;
    10'd26:  neuron_7_mul_25_p <= Pix_726;
    10'd27:  neuron_7_mul_25_p <= Pix_727;
    default: neuron_7_mul_25_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_26_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_26_p <= Pix_728;
    10'd1:  neuron_7_mul_26_p <= Pix_729;
    10'd2:  neuron_7_mul_26_p <= Pix_730;
    10'd3:  neuron_7_mul_26_p <= Pix_731;
    10'd4:  neuron_7_mul_26_p <= Pix_732;
    10'd5:  neuron_7_mul_26_p <= Pix_733;
    10'd6:  neuron_7_mul_26_p <= Pix_734;
    10'd7:  neuron_7_mul_26_p <= Pix_735;
    10'd8:  neuron_7_mul_26_p <= Pix_736;
    10'd9:  neuron_7_mul_26_p <= Pix_737;
    10'd10:  neuron_7_mul_26_p <= Pix_738;
    10'd11:  neuron_7_mul_26_p <= Pix_739;
    10'd12:  neuron_7_mul_26_p <= Pix_740;
    10'd13:  neuron_7_mul_26_p <= Pix_741;
    10'd14:  neuron_7_mul_26_p <= Pix_742;
    10'd15:  neuron_7_mul_26_p <= Pix_743;
    10'd16:  neuron_7_mul_26_p <= Pix_744;
    10'd17:  neuron_7_mul_26_p <= Pix_745;
    10'd18:  neuron_7_mul_26_p <= Pix_746;
    10'd19:  neuron_7_mul_26_p <= Pix_747;
    10'd20:  neuron_7_mul_26_p <= Pix_748;
    10'd21:  neuron_7_mul_26_p <= Pix_749;
    10'd22:  neuron_7_mul_26_p <= Pix_750;
    10'd23:  neuron_7_mul_26_p <= Pix_751;
    10'd24:  neuron_7_mul_26_p <= Pix_752;
    10'd25:  neuron_7_mul_26_p <= Pix_753;
    10'd26:  neuron_7_mul_26_p <= Pix_754;
    10'd27:  neuron_7_mul_26_p <= Pix_755;
    default: neuron_7_mul_26_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_7_mul_27_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_7_mul_27_p <= Pix_756;
    10'd1:  neuron_7_mul_27_p <= Pix_757;
    10'd2:  neuron_7_mul_27_p <= Pix_758;
    10'd3:  neuron_7_mul_27_p <= Pix_759;
    10'd4:  neuron_7_mul_27_p <= Pix_760;
    10'd5:  neuron_7_mul_27_p <= Pix_761;
    10'd6:  neuron_7_mul_27_p <= Pix_762;
    10'd7:  neuron_7_mul_27_p <= Pix_763;
    10'd8:  neuron_7_mul_27_p <= Pix_764;
    10'd9:  neuron_7_mul_27_p <= Pix_765;
    10'd10:  neuron_7_mul_27_p <= Pix_766;
    10'd11:  neuron_7_mul_27_p <= Pix_767;
    10'd12:  neuron_7_mul_27_p <= Pix_768;
    10'd13:  neuron_7_mul_27_p <= Pix_769;
    10'd14:  neuron_7_mul_27_p <= Pix_770;
    10'd15:  neuron_7_mul_27_p <= Pix_771;
    10'd16:  neuron_7_mul_27_p <= Pix_772;
    10'd17:  neuron_7_mul_27_p <= Pix_773;
    10'd18:  neuron_7_mul_27_p <= Pix_774;
    10'd19:  neuron_7_mul_27_p <= Pix_775;
    10'd20:  neuron_7_mul_27_p <= Pix_776;
    10'd21:  neuron_7_mul_27_p <= Pix_777;
    10'd22:  neuron_7_mul_27_p <= Pix_778;
    10'd23:  neuron_7_mul_27_p <= Pix_779;
    10'd24:  neuron_7_mul_27_p <= Pix_780;
    10'd25:  neuron_7_mul_27_p <= Pix_781;
    10'd26:  neuron_7_mul_27_p <= Pix_782;
    10'd27:  neuron_7_mul_27_p <= Pix_783;
    default: neuron_7_mul_27_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_0_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_0_p <= Pix_0;
    10'd1:  neuron_8_mul_0_p <= Pix_1;
    10'd2:  neuron_8_mul_0_p <= Pix_2;
    10'd3:  neuron_8_mul_0_p <= Pix_3;
    10'd4:  neuron_8_mul_0_p <= Pix_4;
    10'd5:  neuron_8_mul_0_p <= Pix_5;
    10'd6:  neuron_8_mul_0_p <= Pix_6;
    10'd7:  neuron_8_mul_0_p <= Pix_7;
    10'd8:  neuron_8_mul_0_p <= Pix_8;
    10'd9:  neuron_8_mul_0_p <= Pix_9;
    10'd10:  neuron_8_mul_0_p <= Pix_10;
    10'd11:  neuron_8_mul_0_p <= Pix_11;
    10'd12:  neuron_8_mul_0_p <= Pix_12;
    10'd13:  neuron_8_mul_0_p <= Pix_13;
    10'd14:  neuron_8_mul_0_p <= Pix_14;
    10'd15:  neuron_8_mul_0_p <= Pix_15;
    10'd16:  neuron_8_mul_0_p <= Pix_16;
    10'd17:  neuron_8_mul_0_p <= Pix_17;
    10'd18:  neuron_8_mul_0_p <= Pix_18;
    10'd19:  neuron_8_mul_0_p <= Pix_19;
    10'd20:  neuron_8_mul_0_p <= Pix_20;
    10'd21:  neuron_8_mul_0_p <= Pix_21;
    10'd22:  neuron_8_mul_0_p <= Pix_22;
    10'd23:  neuron_8_mul_0_p <= Pix_23;
    10'd24:  neuron_8_mul_0_p <= Pix_24;
    10'd25:  neuron_8_mul_0_p <= Pix_25;
    10'd26:  neuron_8_mul_0_p <= Pix_26;
    10'd27:  neuron_8_mul_0_p <= Pix_27;
    default: neuron_8_mul_0_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_1_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_1_p <= Pix_28;
    10'd1:  neuron_8_mul_1_p <= Pix_29;
    10'd2:  neuron_8_mul_1_p <= Pix_30;
    10'd3:  neuron_8_mul_1_p <= Pix_31;
    10'd4:  neuron_8_mul_1_p <= Pix_32;
    10'd5:  neuron_8_mul_1_p <= Pix_33;
    10'd6:  neuron_8_mul_1_p <= Pix_34;
    10'd7:  neuron_8_mul_1_p <= Pix_35;
    10'd8:  neuron_8_mul_1_p <= Pix_36;
    10'd9:  neuron_8_mul_1_p <= Pix_37;
    10'd10:  neuron_8_mul_1_p <= Pix_38;
    10'd11:  neuron_8_mul_1_p <= Pix_39;
    10'd12:  neuron_8_mul_1_p <= Pix_40;
    10'd13:  neuron_8_mul_1_p <= Pix_41;
    10'd14:  neuron_8_mul_1_p <= Pix_42;
    10'd15:  neuron_8_mul_1_p <= Pix_43;
    10'd16:  neuron_8_mul_1_p <= Pix_44;
    10'd17:  neuron_8_mul_1_p <= Pix_45;
    10'd18:  neuron_8_mul_1_p <= Pix_46;
    10'd19:  neuron_8_mul_1_p <= Pix_47;
    10'd20:  neuron_8_mul_1_p <= Pix_48;
    10'd21:  neuron_8_mul_1_p <= Pix_49;
    10'd22:  neuron_8_mul_1_p <= Pix_50;
    10'd23:  neuron_8_mul_1_p <= Pix_51;
    10'd24:  neuron_8_mul_1_p <= Pix_52;
    10'd25:  neuron_8_mul_1_p <= Pix_53;
    10'd26:  neuron_8_mul_1_p <= Pix_54;
    10'd27:  neuron_8_mul_1_p <= Pix_55;
    default: neuron_8_mul_1_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_2_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_2_p <= Pix_56;
    10'd1:  neuron_8_mul_2_p <= Pix_57;
    10'd2:  neuron_8_mul_2_p <= Pix_58;
    10'd3:  neuron_8_mul_2_p <= Pix_59;
    10'd4:  neuron_8_mul_2_p <= Pix_60;
    10'd5:  neuron_8_mul_2_p <= Pix_61;
    10'd6:  neuron_8_mul_2_p <= Pix_62;
    10'd7:  neuron_8_mul_2_p <= Pix_63;
    10'd8:  neuron_8_mul_2_p <= Pix_64;
    10'd9:  neuron_8_mul_2_p <= Pix_65;
    10'd10:  neuron_8_mul_2_p <= Pix_66;
    10'd11:  neuron_8_mul_2_p <= Pix_67;
    10'd12:  neuron_8_mul_2_p <= Pix_68;
    10'd13:  neuron_8_mul_2_p <= Pix_69;
    10'd14:  neuron_8_mul_2_p <= Pix_70;
    10'd15:  neuron_8_mul_2_p <= Pix_71;
    10'd16:  neuron_8_mul_2_p <= Pix_72;
    10'd17:  neuron_8_mul_2_p <= Pix_73;
    10'd18:  neuron_8_mul_2_p <= Pix_74;
    10'd19:  neuron_8_mul_2_p <= Pix_75;
    10'd20:  neuron_8_mul_2_p <= Pix_76;
    10'd21:  neuron_8_mul_2_p <= Pix_77;
    10'd22:  neuron_8_mul_2_p <= Pix_78;
    10'd23:  neuron_8_mul_2_p <= Pix_79;
    10'd24:  neuron_8_mul_2_p <= Pix_80;
    10'd25:  neuron_8_mul_2_p <= Pix_81;
    10'd26:  neuron_8_mul_2_p <= Pix_82;
    10'd27:  neuron_8_mul_2_p <= Pix_83;
    default: neuron_8_mul_2_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_3_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_3_p <= Pix_84;
    10'd1:  neuron_8_mul_3_p <= Pix_85;
    10'd2:  neuron_8_mul_3_p <= Pix_86;
    10'd3:  neuron_8_mul_3_p <= Pix_87;
    10'd4:  neuron_8_mul_3_p <= Pix_88;
    10'd5:  neuron_8_mul_3_p <= Pix_89;
    10'd6:  neuron_8_mul_3_p <= Pix_90;
    10'd7:  neuron_8_mul_3_p <= Pix_91;
    10'd8:  neuron_8_mul_3_p <= Pix_92;
    10'd9:  neuron_8_mul_3_p <= Pix_93;
    10'd10:  neuron_8_mul_3_p <= Pix_94;
    10'd11:  neuron_8_mul_3_p <= Pix_95;
    10'd12:  neuron_8_mul_3_p <= Pix_96;
    10'd13:  neuron_8_mul_3_p <= Pix_97;
    10'd14:  neuron_8_mul_3_p <= Pix_98;
    10'd15:  neuron_8_mul_3_p <= Pix_99;
    10'd16:  neuron_8_mul_3_p <= Pix_100;
    10'd17:  neuron_8_mul_3_p <= Pix_101;
    10'd18:  neuron_8_mul_3_p <= Pix_102;
    10'd19:  neuron_8_mul_3_p <= Pix_103;
    10'd20:  neuron_8_mul_3_p <= Pix_104;
    10'd21:  neuron_8_mul_3_p <= Pix_105;
    10'd22:  neuron_8_mul_3_p <= Pix_106;
    10'd23:  neuron_8_mul_3_p <= Pix_107;
    10'd24:  neuron_8_mul_3_p <= Pix_108;
    10'd25:  neuron_8_mul_3_p <= Pix_109;
    10'd26:  neuron_8_mul_3_p <= Pix_110;
    10'd27:  neuron_8_mul_3_p <= Pix_111;
    default: neuron_8_mul_3_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_4_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_4_p <= Pix_112;
    10'd1:  neuron_8_mul_4_p <= Pix_113;
    10'd2:  neuron_8_mul_4_p <= Pix_114;
    10'd3:  neuron_8_mul_4_p <= Pix_115;
    10'd4:  neuron_8_mul_4_p <= Pix_116;
    10'd5:  neuron_8_mul_4_p <= Pix_117;
    10'd6:  neuron_8_mul_4_p <= Pix_118;
    10'd7:  neuron_8_mul_4_p <= Pix_119;
    10'd8:  neuron_8_mul_4_p <= Pix_120;
    10'd9:  neuron_8_mul_4_p <= Pix_121;
    10'd10:  neuron_8_mul_4_p <= Pix_122;
    10'd11:  neuron_8_mul_4_p <= Pix_123;
    10'd12:  neuron_8_mul_4_p <= Pix_124;
    10'd13:  neuron_8_mul_4_p <= Pix_125;
    10'd14:  neuron_8_mul_4_p <= Pix_126;
    10'd15:  neuron_8_mul_4_p <= Pix_127;
    10'd16:  neuron_8_mul_4_p <= Pix_128;
    10'd17:  neuron_8_mul_4_p <= Pix_129;
    10'd18:  neuron_8_mul_4_p <= Pix_130;
    10'd19:  neuron_8_mul_4_p <= Pix_131;
    10'd20:  neuron_8_mul_4_p <= Pix_132;
    10'd21:  neuron_8_mul_4_p <= Pix_133;
    10'd22:  neuron_8_mul_4_p <= Pix_134;
    10'd23:  neuron_8_mul_4_p <= Pix_135;
    10'd24:  neuron_8_mul_4_p <= Pix_136;
    10'd25:  neuron_8_mul_4_p <= Pix_137;
    10'd26:  neuron_8_mul_4_p <= Pix_138;
    10'd27:  neuron_8_mul_4_p <= Pix_139;
    default: neuron_8_mul_4_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_5_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_5_p <= Pix_140;
    10'd1:  neuron_8_mul_5_p <= Pix_141;
    10'd2:  neuron_8_mul_5_p <= Pix_142;
    10'd3:  neuron_8_mul_5_p <= Pix_143;
    10'd4:  neuron_8_mul_5_p <= Pix_144;
    10'd5:  neuron_8_mul_5_p <= Pix_145;
    10'd6:  neuron_8_mul_5_p <= Pix_146;
    10'd7:  neuron_8_mul_5_p <= Pix_147;
    10'd8:  neuron_8_mul_5_p <= Pix_148;
    10'd9:  neuron_8_mul_5_p <= Pix_149;
    10'd10:  neuron_8_mul_5_p <= Pix_150;
    10'd11:  neuron_8_mul_5_p <= Pix_151;
    10'd12:  neuron_8_mul_5_p <= Pix_152;
    10'd13:  neuron_8_mul_5_p <= Pix_153;
    10'd14:  neuron_8_mul_5_p <= Pix_154;
    10'd15:  neuron_8_mul_5_p <= Pix_155;
    10'd16:  neuron_8_mul_5_p <= Pix_156;
    10'd17:  neuron_8_mul_5_p <= Pix_157;
    10'd18:  neuron_8_mul_5_p <= Pix_158;
    10'd19:  neuron_8_mul_5_p <= Pix_159;
    10'd20:  neuron_8_mul_5_p <= Pix_160;
    10'd21:  neuron_8_mul_5_p <= Pix_161;
    10'd22:  neuron_8_mul_5_p <= Pix_162;
    10'd23:  neuron_8_mul_5_p <= Pix_163;
    10'd24:  neuron_8_mul_5_p <= Pix_164;
    10'd25:  neuron_8_mul_5_p <= Pix_165;
    10'd26:  neuron_8_mul_5_p <= Pix_166;
    10'd27:  neuron_8_mul_5_p <= Pix_167;
    default: neuron_8_mul_5_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_6_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_6_p <= Pix_168;
    10'd1:  neuron_8_mul_6_p <= Pix_169;
    10'd2:  neuron_8_mul_6_p <= Pix_170;
    10'd3:  neuron_8_mul_6_p <= Pix_171;
    10'd4:  neuron_8_mul_6_p <= Pix_172;
    10'd5:  neuron_8_mul_6_p <= Pix_173;
    10'd6:  neuron_8_mul_6_p <= Pix_174;
    10'd7:  neuron_8_mul_6_p <= Pix_175;
    10'd8:  neuron_8_mul_6_p <= Pix_176;
    10'd9:  neuron_8_mul_6_p <= Pix_177;
    10'd10:  neuron_8_mul_6_p <= Pix_178;
    10'd11:  neuron_8_mul_6_p <= Pix_179;
    10'd12:  neuron_8_mul_6_p <= Pix_180;
    10'd13:  neuron_8_mul_6_p <= Pix_181;
    10'd14:  neuron_8_mul_6_p <= Pix_182;
    10'd15:  neuron_8_mul_6_p <= Pix_183;
    10'd16:  neuron_8_mul_6_p <= Pix_184;
    10'd17:  neuron_8_mul_6_p <= Pix_185;
    10'd18:  neuron_8_mul_6_p <= Pix_186;
    10'd19:  neuron_8_mul_6_p <= Pix_187;
    10'd20:  neuron_8_mul_6_p <= Pix_188;
    10'd21:  neuron_8_mul_6_p <= Pix_189;
    10'd22:  neuron_8_mul_6_p <= Pix_190;
    10'd23:  neuron_8_mul_6_p <= Pix_191;
    10'd24:  neuron_8_mul_6_p <= Pix_192;
    10'd25:  neuron_8_mul_6_p <= Pix_193;
    10'd26:  neuron_8_mul_6_p <= Pix_194;
    10'd27:  neuron_8_mul_6_p <= Pix_195;
    default: neuron_8_mul_6_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_7_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_7_p <= Pix_196;
    10'd1:  neuron_8_mul_7_p <= Pix_197;
    10'd2:  neuron_8_mul_7_p <= Pix_198;
    10'd3:  neuron_8_mul_7_p <= Pix_199;
    10'd4:  neuron_8_mul_7_p <= Pix_200;
    10'd5:  neuron_8_mul_7_p <= Pix_201;
    10'd6:  neuron_8_mul_7_p <= Pix_202;
    10'd7:  neuron_8_mul_7_p <= Pix_203;
    10'd8:  neuron_8_mul_7_p <= Pix_204;
    10'd9:  neuron_8_mul_7_p <= Pix_205;
    10'd10:  neuron_8_mul_7_p <= Pix_206;
    10'd11:  neuron_8_mul_7_p <= Pix_207;
    10'd12:  neuron_8_mul_7_p <= Pix_208;
    10'd13:  neuron_8_mul_7_p <= Pix_209;
    10'd14:  neuron_8_mul_7_p <= Pix_210;
    10'd15:  neuron_8_mul_7_p <= Pix_211;
    10'd16:  neuron_8_mul_7_p <= Pix_212;
    10'd17:  neuron_8_mul_7_p <= Pix_213;
    10'd18:  neuron_8_mul_7_p <= Pix_214;
    10'd19:  neuron_8_mul_7_p <= Pix_215;
    10'd20:  neuron_8_mul_7_p <= Pix_216;
    10'd21:  neuron_8_mul_7_p <= Pix_217;
    10'd22:  neuron_8_mul_7_p <= Pix_218;
    10'd23:  neuron_8_mul_7_p <= Pix_219;
    10'd24:  neuron_8_mul_7_p <= Pix_220;
    10'd25:  neuron_8_mul_7_p <= Pix_221;
    10'd26:  neuron_8_mul_7_p <= Pix_222;
    10'd27:  neuron_8_mul_7_p <= Pix_223;
    default: neuron_8_mul_7_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_8_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_8_p <= Pix_224;
    10'd1:  neuron_8_mul_8_p <= Pix_225;
    10'd2:  neuron_8_mul_8_p <= Pix_226;
    10'd3:  neuron_8_mul_8_p <= Pix_227;
    10'd4:  neuron_8_mul_8_p <= Pix_228;
    10'd5:  neuron_8_mul_8_p <= Pix_229;
    10'd6:  neuron_8_mul_8_p <= Pix_230;
    10'd7:  neuron_8_mul_8_p <= Pix_231;
    10'd8:  neuron_8_mul_8_p <= Pix_232;
    10'd9:  neuron_8_mul_8_p <= Pix_233;
    10'd10:  neuron_8_mul_8_p <= Pix_234;
    10'd11:  neuron_8_mul_8_p <= Pix_235;
    10'd12:  neuron_8_mul_8_p <= Pix_236;
    10'd13:  neuron_8_mul_8_p <= Pix_237;
    10'd14:  neuron_8_mul_8_p <= Pix_238;
    10'd15:  neuron_8_mul_8_p <= Pix_239;
    10'd16:  neuron_8_mul_8_p <= Pix_240;
    10'd17:  neuron_8_mul_8_p <= Pix_241;
    10'd18:  neuron_8_mul_8_p <= Pix_242;
    10'd19:  neuron_8_mul_8_p <= Pix_243;
    10'd20:  neuron_8_mul_8_p <= Pix_244;
    10'd21:  neuron_8_mul_8_p <= Pix_245;
    10'd22:  neuron_8_mul_8_p <= Pix_246;
    10'd23:  neuron_8_mul_8_p <= Pix_247;
    10'd24:  neuron_8_mul_8_p <= Pix_248;
    10'd25:  neuron_8_mul_8_p <= Pix_249;
    10'd26:  neuron_8_mul_8_p <= Pix_250;
    10'd27:  neuron_8_mul_8_p <= Pix_251;
    default: neuron_8_mul_8_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_9_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_9_p <= Pix_252;
    10'd1:  neuron_8_mul_9_p <= Pix_253;
    10'd2:  neuron_8_mul_9_p <= Pix_254;
    10'd3:  neuron_8_mul_9_p <= Pix_255;
    10'd4:  neuron_8_mul_9_p <= Pix_256;
    10'd5:  neuron_8_mul_9_p <= Pix_257;
    10'd6:  neuron_8_mul_9_p <= Pix_258;
    10'd7:  neuron_8_mul_9_p <= Pix_259;
    10'd8:  neuron_8_mul_9_p <= Pix_260;
    10'd9:  neuron_8_mul_9_p <= Pix_261;
    10'd10:  neuron_8_mul_9_p <= Pix_262;
    10'd11:  neuron_8_mul_9_p <= Pix_263;
    10'd12:  neuron_8_mul_9_p <= Pix_264;
    10'd13:  neuron_8_mul_9_p <= Pix_265;
    10'd14:  neuron_8_mul_9_p <= Pix_266;
    10'd15:  neuron_8_mul_9_p <= Pix_267;
    10'd16:  neuron_8_mul_9_p <= Pix_268;
    10'd17:  neuron_8_mul_9_p <= Pix_269;
    10'd18:  neuron_8_mul_9_p <= Pix_270;
    10'd19:  neuron_8_mul_9_p <= Pix_271;
    10'd20:  neuron_8_mul_9_p <= Pix_272;
    10'd21:  neuron_8_mul_9_p <= Pix_273;
    10'd22:  neuron_8_mul_9_p <= Pix_274;
    10'd23:  neuron_8_mul_9_p <= Pix_275;
    10'd24:  neuron_8_mul_9_p <= Pix_276;
    10'd25:  neuron_8_mul_9_p <= Pix_277;
    10'd26:  neuron_8_mul_9_p <= Pix_278;
    10'd27:  neuron_8_mul_9_p <= Pix_279;
    default: neuron_8_mul_9_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_10_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_10_p <= Pix_280;
    10'd1:  neuron_8_mul_10_p <= Pix_281;
    10'd2:  neuron_8_mul_10_p <= Pix_282;
    10'd3:  neuron_8_mul_10_p <= Pix_283;
    10'd4:  neuron_8_mul_10_p <= Pix_284;
    10'd5:  neuron_8_mul_10_p <= Pix_285;
    10'd6:  neuron_8_mul_10_p <= Pix_286;
    10'd7:  neuron_8_mul_10_p <= Pix_287;
    10'd8:  neuron_8_mul_10_p <= Pix_288;
    10'd9:  neuron_8_mul_10_p <= Pix_289;
    10'd10:  neuron_8_mul_10_p <= Pix_290;
    10'd11:  neuron_8_mul_10_p <= Pix_291;
    10'd12:  neuron_8_mul_10_p <= Pix_292;
    10'd13:  neuron_8_mul_10_p <= Pix_293;
    10'd14:  neuron_8_mul_10_p <= Pix_294;
    10'd15:  neuron_8_mul_10_p <= Pix_295;
    10'd16:  neuron_8_mul_10_p <= Pix_296;
    10'd17:  neuron_8_mul_10_p <= Pix_297;
    10'd18:  neuron_8_mul_10_p <= Pix_298;
    10'd19:  neuron_8_mul_10_p <= Pix_299;
    10'd20:  neuron_8_mul_10_p <= Pix_300;
    10'd21:  neuron_8_mul_10_p <= Pix_301;
    10'd22:  neuron_8_mul_10_p <= Pix_302;
    10'd23:  neuron_8_mul_10_p <= Pix_303;
    10'd24:  neuron_8_mul_10_p <= Pix_304;
    10'd25:  neuron_8_mul_10_p <= Pix_305;
    10'd26:  neuron_8_mul_10_p <= Pix_306;
    10'd27:  neuron_8_mul_10_p <= Pix_307;
    default: neuron_8_mul_10_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_11_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_11_p <= Pix_308;
    10'd1:  neuron_8_mul_11_p <= Pix_309;
    10'd2:  neuron_8_mul_11_p <= Pix_310;
    10'd3:  neuron_8_mul_11_p <= Pix_311;
    10'd4:  neuron_8_mul_11_p <= Pix_312;
    10'd5:  neuron_8_mul_11_p <= Pix_313;
    10'd6:  neuron_8_mul_11_p <= Pix_314;
    10'd7:  neuron_8_mul_11_p <= Pix_315;
    10'd8:  neuron_8_mul_11_p <= Pix_316;
    10'd9:  neuron_8_mul_11_p <= Pix_317;
    10'd10:  neuron_8_mul_11_p <= Pix_318;
    10'd11:  neuron_8_mul_11_p <= Pix_319;
    10'd12:  neuron_8_mul_11_p <= Pix_320;
    10'd13:  neuron_8_mul_11_p <= Pix_321;
    10'd14:  neuron_8_mul_11_p <= Pix_322;
    10'd15:  neuron_8_mul_11_p <= Pix_323;
    10'd16:  neuron_8_mul_11_p <= Pix_324;
    10'd17:  neuron_8_mul_11_p <= Pix_325;
    10'd18:  neuron_8_mul_11_p <= Pix_326;
    10'd19:  neuron_8_mul_11_p <= Pix_327;
    10'd20:  neuron_8_mul_11_p <= Pix_328;
    10'd21:  neuron_8_mul_11_p <= Pix_329;
    10'd22:  neuron_8_mul_11_p <= Pix_330;
    10'd23:  neuron_8_mul_11_p <= Pix_331;
    10'd24:  neuron_8_mul_11_p <= Pix_332;
    10'd25:  neuron_8_mul_11_p <= Pix_333;
    10'd26:  neuron_8_mul_11_p <= Pix_334;
    10'd27:  neuron_8_mul_11_p <= Pix_335;
    default: neuron_8_mul_11_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_12_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_12_p <= Pix_336;
    10'd1:  neuron_8_mul_12_p <= Pix_337;
    10'd2:  neuron_8_mul_12_p <= Pix_338;
    10'd3:  neuron_8_mul_12_p <= Pix_339;
    10'd4:  neuron_8_mul_12_p <= Pix_340;
    10'd5:  neuron_8_mul_12_p <= Pix_341;
    10'd6:  neuron_8_mul_12_p <= Pix_342;
    10'd7:  neuron_8_mul_12_p <= Pix_343;
    10'd8:  neuron_8_mul_12_p <= Pix_344;
    10'd9:  neuron_8_mul_12_p <= Pix_345;
    10'd10:  neuron_8_mul_12_p <= Pix_346;
    10'd11:  neuron_8_mul_12_p <= Pix_347;
    10'd12:  neuron_8_mul_12_p <= Pix_348;
    10'd13:  neuron_8_mul_12_p <= Pix_349;
    10'd14:  neuron_8_mul_12_p <= Pix_350;
    10'd15:  neuron_8_mul_12_p <= Pix_351;
    10'd16:  neuron_8_mul_12_p <= Pix_352;
    10'd17:  neuron_8_mul_12_p <= Pix_353;
    10'd18:  neuron_8_mul_12_p <= Pix_354;
    10'd19:  neuron_8_mul_12_p <= Pix_355;
    10'd20:  neuron_8_mul_12_p <= Pix_356;
    10'd21:  neuron_8_mul_12_p <= Pix_357;
    10'd22:  neuron_8_mul_12_p <= Pix_358;
    10'd23:  neuron_8_mul_12_p <= Pix_359;
    10'd24:  neuron_8_mul_12_p <= Pix_360;
    10'd25:  neuron_8_mul_12_p <= Pix_361;
    10'd26:  neuron_8_mul_12_p <= Pix_362;
    10'd27:  neuron_8_mul_12_p <= Pix_363;
    default: neuron_8_mul_12_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_13_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_13_p <= Pix_364;
    10'd1:  neuron_8_mul_13_p <= Pix_365;
    10'd2:  neuron_8_mul_13_p <= Pix_366;
    10'd3:  neuron_8_mul_13_p <= Pix_367;
    10'd4:  neuron_8_mul_13_p <= Pix_368;
    10'd5:  neuron_8_mul_13_p <= Pix_369;
    10'd6:  neuron_8_mul_13_p <= Pix_370;
    10'd7:  neuron_8_mul_13_p <= Pix_371;
    10'd8:  neuron_8_mul_13_p <= Pix_372;
    10'd9:  neuron_8_mul_13_p <= Pix_373;
    10'd10:  neuron_8_mul_13_p <= Pix_374;
    10'd11:  neuron_8_mul_13_p <= Pix_375;
    10'd12:  neuron_8_mul_13_p <= Pix_376;
    10'd13:  neuron_8_mul_13_p <= Pix_377;
    10'd14:  neuron_8_mul_13_p <= Pix_378;
    10'd15:  neuron_8_mul_13_p <= Pix_379;
    10'd16:  neuron_8_mul_13_p <= Pix_380;
    10'd17:  neuron_8_mul_13_p <= Pix_381;
    10'd18:  neuron_8_mul_13_p <= Pix_382;
    10'd19:  neuron_8_mul_13_p <= Pix_383;
    10'd20:  neuron_8_mul_13_p <= Pix_384;
    10'd21:  neuron_8_mul_13_p <= Pix_385;
    10'd22:  neuron_8_mul_13_p <= Pix_386;
    10'd23:  neuron_8_mul_13_p <= Pix_387;
    10'd24:  neuron_8_mul_13_p <= Pix_388;
    10'd25:  neuron_8_mul_13_p <= Pix_389;
    10'd26:  neuron_8_mul_13_p <= Pix_390;
    10'd27:  neuron_8_mul_13_p <= Pix_391;
    default: neuron_8_mul_13_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_14_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_14_p <= Pix_392;
    10'd1:  neuron_8_mul_14_p <= Pix_393;
    10'd2:  neuron_8_mul_14_p <= Pix_394;
    10'd3:  neuron_8_mul_14_p <= Pix_395;
    10'd4:  neuron_8_mul_14_p <= Pix_396;
    10'd5:  neuron_8_mul_14_p <= Pix_397;
    10'd6:  neuron_8_mul_14_p <= Pix_398;
    10'd7:  neuron_8_mul_14_p <= Pix_399;
    10'd8:  neuron_8_mul_14_p <= Pix_400;
    10'd9:  neuron_8_mul_14_p <= Pix_401;
    10'd10:  neuron_8_mul_14_p <= Pix_402;
    10'd11:  neuron_8_mul_14_p <= Pix_403;
    10'd12:  neuron_8_mul_14_p <= Pix_404;
    10'd13:  neuron_8_mul_14_p <= Pix_405;
    10'd14:  neuron_8_mul_14_p <= Pix_406;
    10'd15:  neuron_8_mul_14_p <= Pix_407;
    10'd16:  neuron_8_mul_14_p <= Pix_408;
    10'd17:  neuron_8_mul_14_p <= Pix_409;
    10'd18:  neuron_8_mul_14_p <= Pix_410;
    10'd19:  neuron_8_mul_14_p <= Pix_411;
    10'd20:  neuron_8_mul_14_p <= Pix_412;
    10'd21:  neuron_8_mul_14_p <= Pix_413;
    10'd22:  neuron_8_mul_14_p <= Pix_414;
    10'd23:  neuron_8_mul_14_p <= Pix_415;
    10'd24:  neuron_8_mul_14_p <= Pix_416;
    10'd25:  neuron_8_mul_14_p <= Pix_417;
    10'd26:  neuron_8_mul_14_p <= Pix_418;
    10'd27:  neuron_8_mul_14_p <= Pix_419;
    default: neuron_8_mul_14_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_15_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_15_p <= Pix_420;
    10'd1:  neuron_8_mul_15_p <= Pix_421;
    10'd2:  neuron_8_mul_15_p <= Pix_422;
    10'd3:  neuron_8_mul_15_p <= Pix_423;
    10'd4:  neuron_8_mul_15_p <= Pix_424;
    10'd5:  neuron_8_mul_15_p <= Pix_425;
    10'd6:  neuron_8_mul_15_p <= Pix_426;
    10'd7:  neuron_8_mul_15_p <= Pix_427;
    10'd8:  neuron_8_mul_15_p <= Pix_428;
    10'd9:  neuron_8_mul_15_p <= Pix_429;
    10'd10:  neuron_8_mul_15_p <= Pix_430;
    10'd11:  neuron_8_mul_15_p <= Pix_431;
    10'd12:  neuron_8_mul_15_p <= Pix_432;
    10'd13:  neuron_8_mul_15_p <= Pix_433;
    10'd14:  neuron_8_mul_15_p <= Pix_434;
    10'd15:  neuron_8_mul_15_p <= Pix_435;
    10'd16:  neuron_8_mul_15_p <= Pix_436;
    10'd17:  neuron_8_mul_15_p <= Pix_437;
    10'd18:  neuron_8_mul_15_p <= Pix_438;
    10'd19:  neuron_8_mul_15_p <= Pix_439;
    10'd20:  neuron_8_mul_15_p <= Pix_440;
    10'd21:  neuron_8_mul_15_p <= Pix_441;
    10'd22:  neuron_8_mul_15_p <= Pix_442;
    10'd23:  neuron_8_mul_15_p <= Pix_443;
    10'd24:  neuron_8_mul_15_p <= Pix_444;
    10'd25:  neuron_8_mul_15_p <= Pix_445;
    10'd26:  neuron_8_mul_15_p <= Pix_446;
    10'd27:  neuron_8_mul_15_p <= Pix_447;
    default: neuron_8_mul_15_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_16_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_16_p <= Pix_448;
    10'd1:  neuron_8_mul_16_p <= Pix_449;
    10'd2:  neuron_8_mul_16_p <= Pix_450;
    10'd3:  neuron_8_mul_16_p <= Pix_451;
    10'd4:  neuron_8_mul_16_p <= Pix_452;
    10'd5:  neuron_8_mul_16_p <= Pix_453;
    10'd6:  neuron_8_mul_16_p <= Pix_454;
    10'd7:  neuron_8_mul_16_p <= Pix_455;
    10'd8:  neuron_8_mul_16_p <= Pix_456;
    10'd9:  neuron_8_mul_16_p <= Pix_457;
    10'd10:  neuron_8_mul_16_p <= Pix_458;
    10'd11:  neuron_8_mul_16_p <= Pix_459;
    10'd12:  neuron_8_mul_16_p <= Pix_460;
    10'd13:  neuron_8_mul_16_p <= Pix_461;
    10'd14:  neuron_8_mul_16_p <= Pix_462;
    10'd15:  neuron_8_mul_16_p <= Pix_463;
    10'd16:  neuron_8_mul_16_p <= Pix_464;
    10'd17:  neuron_8_mul_16_p <= Pix_465;
    10'd18:  neuron_8_mul_16_p <= Pix_466;
    10'd19:  neuron_8_mul_16_p <= Pix_467;
    10'd20:  neuron_8_mul_16_p <= Pix_468;
    10'd21:  neuron_8_mul_16_p <= Pix_469;
    10'd22:  neuron_8_mul_16_p <= Pix_470;
    10'd23:  neuron_8_mul_16_p <= Pix_471;
    10'd24:  neuron_8_mul_16_p <= Pix_472;
    10'd25:  neuron_8_mul_16_p <= Pix_473;
    10'd26:  neuron_8_mul_16_p <= Pix_474;
    10'd27:  neuron_8_mul_16_p <= Pix_475;
    default: neuron_8_mul_16_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_17_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_17_p <= Pix_476;
    10'd1:  neuron_8_mul_17_p <= Pix_477;
    10'd2:  neuron_8_mul_17_p <= Pix_478;
    10'd3:  neuron_8_mul_17_p <= Pix_479;
    10'd4:  neuron_8_mul_17_p <= Pix_480;
    10'd5:  neuron_8_mul_17_p <= Pix_481;
    10'd6:  neuron_8_mul_17_p <= Pix_482;
    10'd7:  neuron_8_mul_17_p <= Pix_483;
    10'd8:  neuron_8_mul_17_p <= Pix_484;
    10'd9:  neuron_8_mul_17_p <= Pix_485;
    10'd10:  neuron_8_mul_17_p <= Pix_486;
    10'd11:  neuron_8_mul_17_p <= Pix_487;
    10'd12:  neuron_8_mul_17_p <= Pix_488;
    10'd13:  neuron_8_mul_17_p <= Pix_489;
    10'd14:  neuron_8_mul_17_p <= Pix_490;
    10'd15:  neuron_8_mul_17_p <= Pix_491;
    10'd16:  neuron_8_mul_17_p <= Pix_492;
    10'd17:  neuron_8_mul_17_p <= Pix_493;
    10'd18:  neuron_8_mul_17_p <= Pix_494;
    10'd19:  neuron_8_mul_17_p <= Pix_495;
    10'd20:  neuron_8_mul_17_p <= Pix_496;
    10'd21:  neuron_8_mul_17_p <= Pix_497;
    10'd22:  neuron_8_mul_17_p <= Pix_498;
    10'd23:  neuron_8_mul_17_p <= Pix_499;
    10'd24:  neuron_8_mul_17_p <= Pix_500;
    10'd25:  neuron_8_mul_17_p <= Pix_501;
    10'd26:  neuron_8_mul_17_p <= Pix_502;
    10'd27:  neuron_8_mul_17_p <= Pix_503;
    default: neuron_8_mul_17_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_18_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_18_p <= Pix_504;
    10'd1:  neuron_8_mul_18_p <= Pix_505;
    10'd2:  neuron_8_mul_18_p <= Pix_506;
    10'd3:  neuron_8_mul_18_p <= Pix_507;
    10'd4:  neuron_8_mul_18_p <= Pix_508;
    10'd5:  neuron_8_mul_18_p <= Pix_509;
    10'd6:  neuron_8_mul_18_p <= Pix_510;
    10'd7:  neuron_8_mul_18_p <= Pix_511;
    10'd8:  neuron_8_mul_18_p <= Pix_512;
    10'd9:  neuron_8_mul_18_p <= Pix_513;
    10'd10:  neuron_8_mul_18_p <= Pix_514;
    10'd11:  neuron_8_mul_18_p <= Pix_515;
    10'd12:  neuron_8_mul_18_p <= Pix_516;
    10'd13:  neuron_8_mul_18_p <= Pix_517;
    10'd14:  neuron_8_mul_18_p <= Pix_518;
    10'd15:  neuron_8_mul_18_p <= Pix_519;
    10'd16:  neuron_8_mul_18_p <= Pix_520;
    10'd17:  neuron_8_mul_18_p <= Pix_521;
    10'd18:  neuron_8_mul_18_p <= Pix_522;
    10'd19:  neuron_8_mul_18_p <= Pix_523;
    10'd20:  neuron_8_mul_18_p <= Pix_524;
    10'd21:  neuron_8_mul_18_p <= Pix_525;
    10'd22:  neuron_8_mul_18_p <= Pix_526;
    10'd23:  neuron_8_mul_18_p <= Pix_527;
    10'd24:  neuron_8_mul_18_p <= Pix_528;
    10'd25:  neuron_8_mul_18_p <= Pix_529;
    10'd26:  neuron_8_mul_18_p <= Pix_530;
    10'd27:  neuron_8_mul_18_p <= Pix_531;
    default: neuron_8_mul_18_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_19_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_19_p <= Pix_532;
    10'd1:  neuron_8_mul_19_p <= Pix_533;
    10'd2:  neuron_8_mul_19_p <= Pix_534;
    10'd3:  neuron_8_mul_19_p <= Pix_535;
    10'd4:  neuron_8_mul_19_p <= Pix_536;
    10'd5:  neuron_8_mul_19_p <= Pix_537;
    10'd6:  neuron_8_mul_19_p <= Pix_538;
    10'd7:  neuron_8_mul_19_p <= Pix_539;
    10'd8:  neuron_8_mul_19_p <= Pix_540;
    10'd9:  neuron_8_mul_19_p <= Pix_541;
    10'd10:  neuron_8_mul_19_p <= Pix_542;
    10'd11:  neuron_8_mul_19_p <= Pix_543;
    10'd12:  neuron_8_mul_19_p <= Pix_544;
    10'd13:  neuron_8_mul_19_p <= Pix_545;
    10'd14:  neuron_8_mul_19_p <= Pix_546;
    10'd15:  neuron_8_mul_19_p <= Pix_547;
    10'd16:  neuron_8_mul_19_p <= Pix_548;
    10'd17:  neuron_8_mul_19_p <= Pix_549;
    10'd18:  neuron_8_mul_19_p <= Pix_550;
    10'd19:  neuron_8_mul_19_p <= Pix_551;
    10'd20:  neuron_8_mul_19_p <= Pix_552;
    10'd21:  neuron_8_mul_19_p <= Pix_553;
    10'd22:  neuron_8_mul_19_p <= Pix_554;
    10'd23:  neuron_8_mul_19_p <= Pix_555;
    10'd24:  neuron_8_mul_19_p <= Pix_556;
    10'd25:  neuron_8_mul_19_p <= Pix_557;
    10'd26:  neuron_8_mul_19_p <= Pix_558;
    10'd27:  neuron_8_mul_19_p <= Pix_559;
    default: neuron_8_mul_19_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_20_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_20_p <= Pix_560;
    10'd1:  neuron_8_mul_20_p <= Pix_561;
    10'd2:  neuron_8_mul_20_p <= Pix_562;
    10'd3:  neuron_8_mul_20_p <= Pix_563;
    10'd4:  neuron_8_mul_20_p <= Pix_564;
    10'd5:  neuron_8_mul_20_p <= Pix_565;
    10'd6:  neuron_8_mul_20_p <= Pix_566;
    10'd7:  neuron_8_mul_20_p <= Pix_567;
    10'd8:  neuron_8_mul_20_p <= Pix_568;
    10'd9:  neuron_8_mul_20_p <= Pix_569;
    10'd10:  neuron_8_mul_20_p <= Pix_570;
    10'd11:  neuron_8_mul_20_p <= Pix_571;
    10'd12:  neuron_8_mul_20_p <= Pix_572;
    10'd13:  neuron_8_mul_20_p <= Pix_573;
    10'd14:  neuron_8_mul_20_p <= Pix_574;
    10'd15:  neuron_8_mul_20_p <= Pix_575;
    10'd16:  neuron_8_mul_20_p <= Pix_576;
    10'd17:  neuron_8_mul_20_p <= Pix_577;
    10'd18:  neuron_8_mul_20_p <= Pix_578;
    10'd19:  neuron_8_mul_20_p <= Pix_579;
    10'd20:  neuron_8_mul_20_p <= Pix_580;
    10'd21:  neuron_8_mul_20_p <= Pix_581;
    10'd22:  neuron_8_mul_20_p <= Pix_582;
    10'd23:  neuron_8_mul_20_p <= Pix_583;
    10'd24:  neuron_8_mul_20_p <= Pix_584;
    10'd25:  neuron_8_mul_20_p <= Pix_585;
    10'd26:  neuron_8_mul_20_p <= Pix_586;
    10'd27:  neuron_8_mul_20_p <= Pix_587;
    default: neuron_8_mul_20_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_21_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_21_p <= Pix_588;
    10'd1:  neuron_8_mul_21_p <= Pix_589;
    10'd2:  neuron_8_mul_21_p <= Pix_590;
    10'd3:  neuron_8_mul_21_p <= Pix_591;
    10'd4:  neuron_8_mul_21_p <= Pix_592;
    10'd5:  neuron_8_mul_21_p <= Pix_593;
    10'd6:  neuron_8_mul_21_p <= Pix_594;
    10'd7:  neuron_8_mul_21_p <= Pix_595;
    10'd8:  neuron_8_mul_21_p <= Pix_596;
    10'd9:  neuron_8_mul_21_p <= Pix_597;
    10'd10:  neuron_8_mul_21_p <= Pix_598;
    10'd11:  neuron_8_mul_21_p <= Pix_599;
    10'd12:  neuron_8_mul_21_p <= Pix_600;
    10'd13:  neuron_8_mul_21_p <= Pix_601;
    10'd14:  neuron_8_mul_21_p <= Pix_602;
    10'd15:  neuron_8_mul_21_p <= Pix_603;
    10'd16:  neuron_8_mul_21_p <= Pix_604;
    10'd17:  neuron_8_mul_21_p <= Pix_605;
    10'd18:  neuron_8_mul_21_p <= Pix_606;
    10'd19:  neuron_8_mul_21_p <= Pix_607;
    10'd20:  neuron_8_mul_21_p <= Pix_608;
    10'd21:  neuron_8_mul_21_p <= Pix_609;
    10'd22:  neuron_8_mul_21_p <= Pix_610;
    10'd23:  neuron_8_mul_21_p <= Pix_611;
    10'd24:  neuron_8_mul_21_p <= Pix_612;
    10'd25:  neuron_8_mul_21_p <= Pix_613;
    10'd26:  neuron_8_mul_21_p <= Pix_614;
    10'd27:  neuron_8_mul_21_p <= Pix_615;
    default: neuron_8_mul_21_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_22_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_22_p <= Pix_616;
    10'd1:  neuron_8_mul_22_p <= Pix_617;
    10'd2:  neuron_8_mul_22_p <= Pix_618;
    10'd3:  neuron_8_mul_22_p <= Pix_619;
    10'd4:  neuron_8_mul_22_p <= Pix_620;
    10'd5:  neuron_8_mul_22_p <= Pix_621;
    10'd6:  neuron_8_mul_22_p <= Pix_622;
    10'd7:  neuron_8_mul_22_p <= Pix_623;
    10'd8:  neuron_8_mul_22_p <= Pix_624;
    10'd9:  neuron_8_mul_22_p <= Pix_625;
    10'd10:  neuron_8_mul_22_p <= Pix_626;
    10'd11:  neuron_8_mul_22_p <= Pix_627;
    10'd12:  neuron_8_mul_22_p <= Pix_628;
    10'd13:  neuron_8_mul_22_p <= Pix_629;
    10'd14:  neuron_8_mul_22_p <= Pix_630;
    10'd15:  neuron_8_mul_22_p <= Pix_631;
    10'd16:  neuron_8_mul_22_p <= Pix_632;
    10'd17:  neuron_8_mul_22_p <= Pix_633;
    10'd18:  neuron_8_mul_22_p <= Pix_634;
    10'd19:  neuron_8_mul_22_p <= Pix_635;
    10'd20:  neuron_8_mul_22_p <= Pix_636;
    10'd21:  neuron_8_mul_22_p <= Pix_637;
    10'd22:  neuron_8_mul_22_p <= Pix_638;
    10'd23:  neuron_8_mul_22_p <= Pix_639;
    10'd24:  neuron_8_mul_22_p <= Pix_640;
    10'd25:  neuron_8_mul_22_p <= Pix_641;
    10'd26:  neuron_8_mul_22_p <= Pix_642;
    10'd27:  neuron_8_mul_22_p <= Pix_643;
    default: neuron_8_mul_22_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_23_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_23_p <= Pix_644;
    10'd1:  neuron_8_mul_23_p <= Pix_645;
    10'd2:  neuron_8_mul_23_p <= Pix_646;
    10'd3:  neuron_8_mul_23_p <= Pix_647;
    10'd4:  neuron_8_mul_23_p <= Pix_648;
    10'd5:  neuron_8_mul_23_p <= Pix_649;
    10'd6:  neuron_8_mul_23_p <= Pix_650;
    10'd7:  neuron_8_mul_23_p <= Pix_651;
    10'd8:  neuron_8_mul_23_p <= Pix_652;
    10'd9:  neuron_8_mul_23_p <= Pix_653;
    10'd10:  neuron_8_mul_23_p <= Pix_654;
    10'd11:  neuron_8_mul_23_p <= Pix_655;
    10'd12:  neuron_8_mul_23_p <= Pix_656;
    10'd13:  neuron_8_mul_23_p <= Pix_657;
    10'd14:  neuron_8_mul_23_p <= Pix_658;
    10'd15:  neuron_8_mul_23_p <= Pix_659;
    10'd16:  neuron_8_mul_23_p <= Pix_660;
    10'd17:  neuron_8_mul_23_p <= Pix_661;
    10'd18:  neuron_8_mul_23_p <= Pix_662;
    10'd19:  neuron_8_mul_23_p <= Pix_663;
    10'd20:  neuron_8_mul_23_p <= Pix_664;
    10'd21:  neuron_8_mul_23_p <= Pix_665;
    10'd22:  neuron_8_mul_23_p <= Pix_666;
    10'd23:  neuron_8_mul_23_p <= Pix_667;
    10'd24:  neuron_8_mul_23_p <= Pix_668;
    10'd25:  neuron_8_mul_23_p <= Pix_669;
    10'd26:  neuron_8_mul_23_p <= Pix_670;
    10'd27:  neuron_8_mul_23_p <= Pix_671;
    default: neuron_8_mul_23_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_24_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_24_p <= Pix_672;
    10'd1:  neuron_8_mul_24_p <= Pix_673;
    10'd2:  neuron_8_mul_24_p <= Pix_674;
    10'd3:  neuron_8_mul_24_p <= Pix_675;
    10'd4:  neuron_8_mul_24_p <= Pix_676;
    10'd5:  neuron_8_mul_24_p <= Pix_677;
    10'd6:  neuron_8_mul_24_p <= Pix_678;
    10'd7:  neuron_8_mul_24_p <= Pix_679;
    10'd8:  neuron_8_mul_24_p <= Pix_680;
    10'd9:  neuron_8_mul_24_p <= Pix_681;
    10'd10:  neuron_8_mul_24_p <= Pix_682;
    10'd11:  neuron_8_mul_24_p <= Pix_683;
    10'd12:  neuron_8_mul_24_p <= Pix_684;
    10'd13:  neuron_8_mul_24_p <= Pix_685;
    10'd14:  neuron_8_mul_24_p <= Pix_686;
    10'd15:  neuron_8_mul_24_p <= Pix_687;
    10'd16:  neuron_8_mul_24_p <= Pix_688;
    10'd17:  neuron_8_mul_24_p <= Pix_689;
    10'd18:  neuron_8_mul_24_p <= Pix_690;
    10'd19:  neuron_8_mul_24_p <= Pix_691;
    10'd20:  neuron_8_mul_24_p <= Pix_692;
    10'd21:  neuron_8_mul_24_p <= Pix_693;
    10'd22:  neuron_8_mul_24_p <= Pix_694;
    10'd23:  neuron_8_mul_24_p <= Pix_695;
    10'd24:  neuron_8_mul_24_p <= Pix_696;
    10'd25:  neuron_8_mul_24_p <= Pix_697;
    10'd26:  neuron_8_mul_24_p <= Pix_698;
    10'd27:  neuron_8_mul_24_p <= Pix_699;
    default: neuron_8_mul_24_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_25_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_25_p <= Pix_700;
    10'd1:  neuron_8_mul_25_p <= Pix_701;
    10'd2:  neuron_8_mul_25_p <= Pix_702;
    10'd3:  neuron_8_mul_25_p <= Pix_703;
    10'd4:  neuron_8_mul_25_p <= Pix_704;
    10'd5:  neuron_8_mul_25_p <= Pix_705;
    10'd6:  neuron_8_mul_25_p <= Pix_706;
    10'd7:  neuron_8_mul_25_p <= Pix_707;
    10'd8:  neuron_8_mul_25_p <= Pix_708;
    10'd9:  neuron_8_mul_25_p <= Pix_709;
    10'd10:  neuron_8_mul_25_p <= Pix_710;
    10'd11:  neuron_8_mul_25_p <= Pix_711;
    10'd12:  neuron_8_mul_25_p <= Pix_712;
    10'd13:  neuron_8_mul_25_p <= Pix_713;
    10'd14:  neuron_8_mul_25_p <= Pix_714;
    10'd15:  neuron_8_mul_25_p <= Pix_715;
    10'd16:  neuron_8_mul_25_p <= Pix_716;
    10'd17:  neuron_8_mul_25_p <= Pix_717;
    10'd18:  neuron_8_mul_25_p <= Pix_718;
    10'd19:  neuron_8_mul_25_p <= Pix_719;
    10'd20:  neuron_8_mul_25_p <= Pix_720;
    10'd21:  neuron_8_mul_25_p <= Pix_721;
    10'd22:  neuron_8_mul_25_p <= Pix_722;
    10'd23:  neuron_8_mul_25_p <= Pix_723;
    10'd24:  neuron_8_mul_25_p <= Pix_724;
    10'd25:  neuron_8_mul_25_p <= Pix_725;
    10'd26:  neuron_8_mul_25_p <= Pix_726;
    10'd27:  neuron_8_mul_25_p <= Pix_727;
    default: neuron_8_mul_25_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_26_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_26_p <= Pix_728;
    10'd1:  neuron_8_mul_26_p <= Pix_729;
    10'd2:  neuron_8_mul_26_p <= Pix_730;
    10'd3:  neuron_8_mul_26_p <= Pix_731;
    10'd4:  neuron_8_mul_26_p <= Pix_732;
    10'd5:  neuron_8_mul_26_p <= Pix_733;
    10'd6:  neuron_8_mul_26_p <= Pix_734;
    10'd7:  neuron_8_mul_26_p <= Pix_735;
    10'd8:  neuron_8_mul_26_p <= Pix_736;
    10'd9:  neuron_8_mul_26_p <= Pix_737;
    10'd10:  neuron_8_mul_26_p <= Pix_738;
    10'd11:  neuron_8_mul_26_p <= Pix_739;
    10'd12:  neuron_8_mul_26_p <= Pix_740;
    10'd13:  neuron_8_mul_26_p <= Pix_741;
    10'd14:  neuron_8_mul_26_p <= Pix_742;
    10'd15:  neuron_8_mul_26_p <= Pix_743;
    10'd16:  neuron_8_mul_26_p <= Pix_744;
    10'd17:  neuron_8_mul_26_p <= Pix_745;
    10'd18:  neuron_8_mul_26_p <= Pix_746;
    10'd19:  neuron_8_mul_26_p <= Pix_747;
    10'd20:  neuron_8_mul_26_p <= Pix_748;
    10'd21:  neuron_8_mul_26_p <= Pix_749;
    10'd22:  neuron_8_mul_26_p <= Pix_750;
    10'd23:  neuron_8_mul_26_p <= Pix_751;
    10'd24:  neuron_8_mul_26_p <= Pix_752;
    10'd25:  neuron_8_mul_26_p <= Pix_753;
    10'd26:  neuron_8_mul_26_p <= Pix_754;
    10'd27:  neuron_8_mul_26_p <= Pix_755;
    default: neuron_8_mul_26_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_8_mul_27_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_8_mul_27_p <= Pix_756;
    10'd1:  neuron_8_mul_27_p <= Pix_757;
    10'd2:  neuron_8_mul_27_p <= Pix_758;
    10'd3:  neuron_8_mul_27_p <= Pix_759;
    10'd4:  neuron_8_mul_27_p <= Pix_760;
    10'd5:  neuron_8_mul_27_p <= Pix_761;
    10'd6:  neuron_8_mul_27_p <= Pix_762;
    10'd7:  neuron_8_mul_27_p <= Pix_763;
    10'd8:  neuron_8_mul_27_p <= Pix_764;
    10'd9:  neuron_8_mul_27_p <= Pix_765;
    10'd10:  neuron_8_mul_27_p <= Pix_766;
    10'd11:  neuron_8_mul_27_p <= Pix_767;
    10'd12:  neuron_8_mul_27_p <= Pix_768;
    10'd13:  neuron_8_mul_27_p <= Pix_769;
    10'd14:  neuron_8_mul_27_p <= Pix_770;
    10'd15:  neuron_8_mul_27_p <= Pix_771;
    10'd16:  neuron_8_mul_27_p <= Pix_772;
    10'd17:  neuron_8_mul_27_p <= Pix_773;
    10'd18:  neuron_8_mul_27_p <= Pix_774;
    10'd19:  neuron_8_mul_27_p <= Pix_775;
    10'd20:  neuron_8_mul_27_p <= Pix_776;
    10'd21:  neuron_8_mul_27_p <= Pix_777;
    10'd22:  neuron_8_mul_27_p <= Pix_778;
    10'd23:  neuron_8_mul_27_p <= Pix_779;
    10'd24:  neuron_8_mul_27_p <= Pix_780;
    10'd25:  neuron_8_mul_27_p <= Pix_781;
    10'd26:  neuron_8_mul_27_p <= Pix_782;
    10'd27:  neuron_8_mul_27_p <= Pix_783;
    default: neuron_8_mul_27_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_0_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_0_p <= Pix_0;
    10'd1:  neuron_9_mul_0_p <= Pix_1;
    10'd2:  neuron_9_mul_0_p <= Pix_2;
    10'd3:  neuron_9_mul_0_p <= Pix_3;
    10'd4:  neuron_9_mul_0_p <= Pix_4;
    10'd5:  neuron_9_mul_0_p <= Pix_5;
    10'd6:  neuron_9_mul_0_p <= Pix_6;
    10'd7:  neuron_9_mul_0_p <= Pix_7;
    10'd8:  neuron_9_mul_0_p <= Pix_8;
    10'd9:  neuron_9_mul_0_p <= Pix_9;
    10'd10:  neuron_9_mul_0_p <= Pix_10;
    10'd11:  neuron_9_mul_0_p <= Pix_11;
    10'd12:  neuron_9_mul_0_p <= Pix_12;
    10'd13:  neuron_9_mul_0_p <= Pix_13;
    10'd14:  neuron_9_mul_0_p <= Pix_14;
    10'd15:  neuron_9_mul_0_p <= Pix_15;
    10'd16:  neuron_9_mul_0_p <= Pix_16;
    10'd17:  neuron_9_mul_0_p <= Pix_17;
    10'd18:  neuron_9_mul_0_p <= Pix_18;
    10'd19:  neuron_9_mul_0_p <= Pix_19;
    10'd20:  neuron_9_mul_0_p <= Pix_20;
    10'd21:  neuron_9_mul_0_p <= Pix_21;
    10'd22:  neuron_9_mul_0_p <= Pix_22;
    10'd23:  neuron_9_mul_0_p <= Pix_23;
    10'd24:  neuron_9_mul_0_p <= Pix_24;
    10'd25:  neuron_9_mul_0_p <= Pix_25;
    10'd26:  neuron_9_mul_0_p <= Pix_26;
    10'd27:  neuron_9_mul_0_p <= Pix_27;
    default: neuron_9_mul_0_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_1_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_1_p <= Pix_28;
    10'd1:  neuron_9_mul_1_p <= Pix_29;
    10'd2:  neuron_9_mul_1_p <= Pix_30;
    10'd3:  neuron_9_mul_1_p <= Pix_31;
    10'd4:  neuron_9_mul_1_p <= Pix_32;
    10'd5:  neuron_9_mul_1_p <= Pix_33;
    10'd6:  neuron_9_mul_1_p <= Pix_34;
    10'd7:  neuron_9_mul_1_p <= Pix_35;
    10'd8:  neuron_9_mul_1_p <= Pix_36;
    10'd9:  neuron_9_mul_1_p <= Pix_37;
    10'd10:  neuron_9_mul_1_p <= Pix_38;
    10'd11:  neuron_9_mul_1_p <= Pix_39;
    10'd12:  neuron_9_mul_1_p <= Pix_40;
    10'd13:  neuron_9_mul_1_p <= Pix_41;
    10'd14:  neuron_9_mul_1_p <= Pix_42;
    10'd15:  neuron_9_mul_1_p <= Pix_43;
    10'd16:  neuron_9_mul_1_p <= Pix_44;
    10'd17:  neuron_9_mul_1_p <= Pix_45;
    10'd18:  neuron_9_mul_1_p <= Pix_46;
    10'd19:  neuron_9_mul_1_p <= Pix_47;
    10'd20:  neuron_9_mul_1_p <= Pix_48;
    10'd21:  neuron_9_mul_1_p <= Pix_49;
    10'd22:  neuron_9_mul_1_p <= Pix_50;
    10'd23:  neuron_9_mul_1_p <= Pix_51;
    10'd24:  neuron_9_mul_1_p <= Pix_52;
    10'd25:  neuron_9_mul_1_p <= Pix_53;
    10'd26:  neuron_9_mul_1_p <= Pix_54;
    10'd27:  neuron_9_mul_1_p <= Pix_55;
    default: neuron_9_mul_1_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_2_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_2_p <= Pix_56;
    10'd1:  neuron_9_mul_2_p <= Pix_57;
    10'd2:  neuron_9_mul_2_p <= Pix_58;
    10'd3:  neuron_9_mul_2_p <= Pix_59;
    10'd4:  neuron_9_mul_2_p <= Pix_60;
    10'd5:  neuron_9_mul_2_p <= Pix_61;
    10'd6:  neuron_9_mul_2_p <= Pix_62;
    10'd7:  neuron_9_mul_2_p <= Pix_63;
    10'd8:  neuron_9_mul_2_p <= Pix_64;
    10'd9:  neuron_9_mul_2_p <= Pix_65;
    10'd10:  neuron_9_mul_2_p <= Pix_66;
    10'd11:  neuron_9_mul_2_p <= Pix_67;
    10'd12:  neuron_9_mul_2_p <= Pix_68;
    10'd13:  neuron_9_mul_2_p <= Pix_69;
    10'd14:  neuron_9_mul_2_p <= Pix_70;
    10'd15:  neuron_9_mul_2_p <= Pix_71;
    10'd16:  neuron_9_mul_2_p <= Pix_72;
    10'd17:  neuron_9_mul_2_p <= Pix_73;
    10'd18:  neuron_9_mul_2_p <= Pix_74;
    10'd19:  neuron_9_mul_2_p <= Pix_75;
    10'd20:  neuron_9_mul_2_p <= Pix_76;
    10'd21:  neuron_9_mul_2_p <= Pix_77;
    10'd22:  neuron_9_mul_2_p <= Pix_78;
    10'd23:  neuron_9_mul_2_p <= Pix_79;
    10'd24:  neuron_9_mul_2_p <= Pix_80;
    10'd25:  neuron_9_mul_2_p <= Pix_81;
    10'd26:  neuron_9_mul_2_p <= Pix_82;
    10'd27:  neuron_9_mul_2_p <= Pix_83;
    default: neuron_9_mul_2_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_3_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_3_p <= Pix_84;
    10'd1:  neuron_9_mul_3_p <= Pix_85;
    10'd2:  neuron_9_mul_3_p <= Pix_86;
    10'd3:  neuron_9_mul_3_p <= Pix_87;
    10'd4:  neuron_9_mul_3_p <= Pix_88;
    10'd5:  neuron_9_mul_3_p <= Pix_89;
    10'd6:  neuron_9_mul_3_p <= Pix_90;
    10'd7:  neuron_9_mul_3_p <= Pix_91;
    10'd8:  neuron_9_mul_3_p <= Pix_92;
    10'd9:  neuron_9_mul_3_p <= Pix_93;
    10'd10:  neuron_9_mul_3_p <= Pix_94;
    10'd11:  neuron_9_mul_3_p <= Pix_95;
    10'd12:  neuron_9_mul_3_p <= Pix_96;
    10'd13:  neuron_9_mul_3_p <= Pix_97;
    10'd14:  neuron_9_mul_3_p <= Pix_98;
    10'd15:  neuron_9_mul_3_p <= Pix_99;
    10'd16:  neuron_9_mul_3_p <= Pix_100;
    10'd17:  neuron_9_mul_3_p <= Pix_101;
    10'd18:  neuron_9_mul_3_p <= Pix_102;
    10'd19:  neuron_9_mul_3_p <= Pix_103;
    10'd20:  neuron_9_mul_3_p <= Pix_104;
    10'd21:  neuron_9_mul_3_p <= Pix_105;
    10'd22:  neuron_9_mul_3_p <= Pix_106;
    10'd23:  neuron_9_mul_3_p <= Pix_107;
    10'd24:  neuron_9_mul_3_p <= Pix_108;
    10'd25:  neuron_9_mul_3_p <= Pix_109;
    10'd26:  neuron_9_mul_3_p <= Pix_110;
    10'd27:  neuron_9_mul_3_p <= Pix_111;
    default: neuron_9_mul_3_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_4_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_4_p <= Pix_112;
    10'd1:  neuron_9_mul_4_p <= Pix_113;
    10'd2:  neuron_9_mul_4_p <= Pix_114;
    10'd3:  neuron_9_mul_4_p <= Pix_115;
    10'd4:  neuron_9_mul_4_p <= Pix_116;
    10'd5:  neuron_9_mul_4_p <= Pix_117;
    10'd6:  neuron_9_mul_4_p <= Pix_118;
    10'd7:  neuron_9_mul_4_p <= Pix_119;
    10'd8:  neuron_9_mul_4_p <= Pix_120;
    10'd9:  neuron_9_mul_4_p <= Pix_121;
    10'd10:  neuron_9_mul_4_p <= Pix_122;
    10'd11:  neuron_9_mul_4_p <= Pix_123;
    10'd12:  neuron_9_mul_4_p <= Pix_124;
    10'd13:  neuron_9_mul_4_p <= Pix_125;
    10'd14:  neuron_9_mul_4_p <= Pix_126;
    10'd15:  neuron_9_mul_4_p <= Pix_127;
    10'd16:  neuron_9_mul_4_p <= Pix_128;
    10'd17:  neuron_9_mul_4_p <= Pix_129;
    10'd18:  neuron_9_mul_4_p <= Pix_130;
    10'd19:  neuron_9_mul_4_p <= Pix_131;
    10'd20:  neuron_9_mul_4_p <= Pix_132;
    10'd21:  neuron_9_mul_4_p <= Pix_133;
    10'd22:  neuron_9_mul_4_p <= Pix_134;
    10'd23:  neuron_9_mul_4_p <= Pix_135;
    10'd24:  neuron_9_mul_4_p <= Pix_136;
    10'd25:  neuron_9_mul_4_p <= Pix_137;
    10'd26:  neuron_9_mul_4_p <= Pix_138;
    10'd27:  neuron_9_mul_4_p <= Pix_139;
    default: neuron_9_mul_4_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_5_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_5_p <= Pix_140;
    10'd1:  neuron_9_mul_5_p <= Pix_141;
    10'd2:  neuron_9_mul_5_p <= Pix_142;
    10'd3:  neuron_9_mul_5_p <= Pix_143;
    10'd4:  neuron_9_mul_5_p <= Pix_144;
    10'd5:  neuron_9_mul_5_p <= Pix_145;
    10'd6:  neuron_9_mul_5_p <= Pix_146;
    10'd7:  neuron_9_mul_5_p <= Pix_147;
    10'd8:  neuron_9_mul_5_p <= Pix_148;
    10'd9:  neuron_9_mul_5_p <= Pix_149;
    10'd10:  neuron_9_mul_5_p <= Pix_150;
    10'd11:  neuron_9_mul_5_p <= Pix_151;
    10'd12:  neuron_9_mul_5_p <= Pix_152;
    10'd13:  neuron_9_mul_5_p <= Pix_153;
    10'd14:  neuron_9_mul_5_p <= Pix_154;
    10'd15:  neuron_9_mul_5_p <= Pix_155;
    10'd16:  neuron_9_mul_5_p <= Pix_156;
    10'd17:  neuron_9_mul_5_p <= Pix_157;
    10'd18:  neuron_9_mul_5_p <= Pix_158;
    10'd19:  neuron_9_mul_5_p <= Pix_159;
    10'd20:  neuron_9_mul_5_p <= Pix_160;
    10'd21:  neuron_9_mul_5_p <= Pix_161;
    10'd22:  neuron_9_mul_5_p <= Pix_162;
    10'd23:  neuron_9_mul_5_p <= Pix_163;
    10'd24:  neuron_9_mul_5_p <= Pix_164;
    10'd25:  neuron_9_mul_5_p <= Pix_165;
    10'd26:  neuron_9_mul_5_p <= Pix_166;
    10'd27:  neuron_9_mul_5_p <= Pix_167;
    default: neuron_9_mul_5_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_6_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_6_p <= Pix_168;
    10'd1:  neuron_9_mul_6_p <= Pix_169;
    10'd2:  neuron_9_mul_6_p <= Pix_170;
    10'd3:  neuron_9_mul_6_p <= Pix_171;
    10'd4:  neuron_9_mul_6_p <= Pix_172;
    10'd5:  neuron_9_mul_6_p <= Pix_173;
    10'd6:  neuron_9_mul_6_p <= Pix_174;
    10'd7:  neuron_9_mul_6_p <= Pix_175;
    10'd8:  neuron_9_mul_6_p <= Pix_176;
    10'd9:  neuron_9_mul_6_p <= Pix_177;
    10'd10:  neuron_9_mul_6_p <= Pix_178;
    10'd11:  neuron_9_mul_6_p <= Pix_179;
    10'd12:  neuron_9_mul_6_p <= Pix_180;
    10'd13:  neuron_9_mul_6_p <= Pix_181;
    10'd14:  neuron_9_mul_6_p <= Pix_182;
    10'd15:  neuron_9_mul_6_p <= Pix_183;
    10'd16:  neuron_9_mul_6_p <= Pix_184;
    10'd17:  neuron_9_mul_6_p <= Pix_185;
    10'd18:  neuron_9_mul_6_p <= Pix_186;
    10'd19:  neuron_9_mul_6_p <= Pix_187;
    10'd20:  neuron_9_mul_6_p <= Pix_188;
    10'd21:  neuron_9_mul_6_p <= Pix_189;
    10'd22:  neuron_9_mul_6_p <= Pix_190;
    10'd23:  neuron_9_mul_6_p <= Pix_191;
    10'd24:  neuron_9_mul_6_p <= Pix_192;
    10'd25:  neuron_9_mul_6_p <= Pix_193;
    10'd26:  neuron_9_mul_6_p <= Pix_194;
    10'd27:  neuron_9_mul_6_p <= Pix_195;
    default: neuron_9_mul_6_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_7_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_7_p <= Pix_196;
    10'd1:  neuron_9_mul_7_p <= Pix_197;
    10'd2:  neuron_9_mul_7_p <= Pix_198;
    10'd3:  neuron_9_mul_7_p <= Pix_199;
    10'd4:  neuron_9_mul_7_p <= Pix_200;
    10'd5:  neuron_9_mul_7_p <= Pix_201;
    10'd6:  neuron_9_mul_7_p <= Pix_202;
    10'd7:  neuron_9_mul_7_p <= Pix_203;
    10'd8:  neuron_9_mul_7_p <= Pix_204;
    10'd9:  neuron_9_mul_7_p <= Pix_205;
    10'd10:  neuron_9_mul_7_p <= Pix_206;
    10'd11:  neuron_9_mul_7_p <= Pix_207;
    10'd12:  neuron_9_mul_7_p <= Pix_208;
    10'd13:  neuron_9_mul_7_p <= Pix_209;
    10'd14:  neuron_9_mul_7_p <= Pix_210;
    10'd15:  neuron_9_mul_7_p <= Pix_211;
    10'd16:  neuron_9_mul_7_p <= Pix_212;
    10'd17:  neuron_9_mul_7_p <= Pix_213;
    10'd18:  neuron_9_mul_7_p <= Pix_214;
    10'd19:  neuron_9_mul_7_p <= Pix_215;
    10'd20:  neuron_9_mul_7_p <= Pix_216;
    10'd21:  neuron_9_mul_7_p <= Pix_217;
    10'd22:  neuron_9_mul_7_p <= Pix_218;
    10'd23:  neuron_9_mul_7_p <= Pix_219;
    10'd24:  neuron_9_mul_7_p <= Pix_220;
    10'd25:  neuron_9_mul_7_p <= Pix_221;
    10'd26:  neuron_9_mul_7_p <= Pix_222;
    10'd27:  neuron_9_mul_7_p <= Pix_223;
    default: neuron_9_mul_7_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_8_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_8_p <= Pix_224;
    10'd1:  neuron_9_mul_8_p <= Pix_225;
    10'd2:  neuron_9_mul_8_p <= Pix_226;
    10'd3:  neuron_9_mul_8_p <= Pix_227;
    10'd4:  neuron_9_mul_8_p <= Pix_228;
    10'd5:  neuron_9_mul_8_p <= Pix_229;
    10'd6:  neuron_9_mul_8_p <= Pix_230;
    10'd7:  neuron_9_mul_8_p <= Pix_231;
    10'd8:  neuron_9_mul_8_p <= Pix_232;
    10'd9:  neuron_9_mul_8_p <= Pix_233;
    10'd10:  neuron_9_mul_8_p <= Pix_234;
    10'd11:  neuron_9_mul_8_p <= Pix_235;
    10'd12:  neuron_9_mul_8_p <= Pix_236;
    10'd13:  neuron_9_mul_8_p <= Pix_237;
    10'd14:  neuron_9_mul_8_p <= Pix_238;
    10'd15:  neuron_9_mul_8_p <= Pix_239;
    10'd16:  neuron_9_mul_8_p <= Pix_240;
    10'd17:  neuron_9_mul_8_p <= Pix_241;
    10'd18:  neuron_9_mul_8_p <= Pix_242;
    10'd19:  neuron_9_mul_8_p <= Pix_243;
    10'd20:  neuron_9_mul_8_p <= Pix_244;
    10'd21:  neuron_9_mul_8_p <= Pix_245;
    10'd22:  neuron_9_mul_8_p <= Pix_246;
    10'd23:  neuron_9_mul_8_p <= Pix_247;
    10'd24:  neuron_9_mul_8_p <= Pix_248;
    10'd25:  neuron_9_mul_8_p <= Pix_249;
    10'd26:  neuron_9_mul_8_p <= Pix_250;
    10'd27:  neuron_9_mul_8_p <= Pix_251;
    default: neuron_9_mul_8_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_9_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_9_p <= Pix_252;
    10'd1:  neuron_9_mul_9_p <= Pix_253;
    10'd2:  neuron_9_mul_9_p <= Pix_254;
    10'd3:  neuron_9_mul_9_p <= Pix_255;
    10'd4:  neuron_9_mul_9_p <= Pix_256;
    10'd5:  neuron_9_mul_9_p <= Pix_257;
    10'd6:  neuron_9_mul_9_p <= Pix_258;
    10'd7:  neuron_9_mul_9_p <= Pix_259;
    10'd8:  neuron_9_mul_9_p <= Pix_260;
    10'd9:  neuron_9_mul_9_p <= Pix_261;
    10'd10:  neuron_9_mul_9_p <= Pix_262;
    10'd11:  neuron_9_mul_9_p <= Pix_263;
    10'd12:  neuron_9_mul_9_p <= Pix_264;
    10'd13:  neuron_9_mul_9_p <= Pix_265;
    10'd14:  neuron_9_mul_9_p <= Pix_266;
    10'd15:  neuron_9_mul_9_p <= Pix_267;
    10'd16:  neuron_9_mul_9_p <= Pix_268;
    10'd17:  neuron_9_mul_9_p <= Pix_269;
    10'd18:  neuron_9_mul_9_p <= Pix_270;
    10'd19:  neuron_9_mul_9_p <= Pix_271;
    10'd20:  neuron_9_mul_9_p <= Pix_272;
    10'd21:  neuron_9_mul_9_p <= Pix_273;
    10'd22:  neuron_9_mul_9_p <= Pix_274;
    10'd23:  neuron_9_mul_9_p <= Pix_275;
    10'd24:  neuron_9_mul_9_p <= Pix_276;
    10'd25:  neuron_9_mul_9_p <= Pix_277;
    10'd26:  neuron_9_mul_9_p <= Pix_278;
    10'd27:  neuron_9_mul_9_p <= Pix_279;
    default: neuron_9_mul_9_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_10_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_10_p <= Pix_280;
    10'd1:  neuron_9_mul_10_p <= Pix_281;
    10'd2:  neuron_9_mul_10_p <= Pix_282;
    10'd3:  neuron_9_mul_10_p <= Pix_283;
    10'd4:  neuron_9_mul_10_p <= Pix_284;
    10'd5:  neuron_9_mul_10_p <= Pix_285;
    10'd6:  neuron_9_mul_10_p <= Pix_286;
    10'd7:  neuron_9_mul_10_p <= Pix_287;
    10'd8:  neuron_9_mul_10_p <= Pix_288;
    10'd9:  neuron_9_mul_10_p <= Pix_289;
    10'd10:  neuron_9_mul_10_p <= Pix_290;
    10'd11:  neuron_9_mul_10_p <= Pix_291;
    10'd12:  neuron_9_mul_10_p <= Pix_292;
    10'd13:  neuron_9_mul_10_p <= Pix_293;
    10'd14:  neuron_9_mul_10_p <= Pix_294;
    10'd15:  neuron_9_mul_10_p <= Pix_295;
    10'd16:  neuron_9_mul_10_p <= Pix_296;
    10'd17:  neuron_9_mul_10_p <= Pix_297;
    10'd18:  neuron_9_mul_10_p <= Pix_298;
    10'd19:  neuron_9_mul_10_p <= Pix_299;
    10'd20:  neuron_9_mul_10_p <= Pix_300;
    10'd21:  neuron_9_mul_10_p <= Pix_301;
    10'd22:  neuron_9_mul_10_p <= Pix_302;
    10'd23:  neuron_9_mul_10_p <= Pix_303;
    10'd24:  neuron_9_mul_10_p <= Pix_304;
    10'd25:  neuron_9_mul_10_p <= Pix_305;
    10'd26:  neuron_9_mul_10_p <= Pix_306;
    10'd27:  neuron_9_mul_10_p <= Pix_307;
    default: neuron_9_mul_10_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_11_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_11_p <= Pix_308;
    10'd1:  neuron_9_mul_11_p <= Pix_309;
    10'd2:  neuron_9_mul_11_p <= Pix_310;
    10'd3:  neuron_9_mul_11_p <= Pix_311;
    10'd4:  neuron_9_mul_11_p <= Pix_312;
    10'd5:  neuron_9_mul_11_p <= Pix_313;
    10'd6:  neuron_9_mul_11_p <= Pix_314;
    10'd7:  neuron_9_mul_11_p <= Pix_315;
    10'd8:  neuron_9_mul_11_p <= Pix_316;
    10'd9:  neuron_9_mul_11_p <= Pix_317;
    10'd10:  neuron_9_mul_11_p <= Pix_318;
    10'd11:  neuron_9_mul_11_p <= Pix_319;
    10'd12:  neuron_9_mul_11_p <= Pix_320;
    10'd13:  neuron_9_mul_11_p <= Pix_321;
    10'd14:  neuron_9_mul_11_p <= Pix_322;
    10'd15:  neuron_9_mul_11_p <= Pix_323;
    10'd16:  neuron_9_mul_11_p <= Pix_324;
    10'd17:  neuron_9_mul_11_p <= Pix_325;
    10'd18:  neuron_9_mul_11_p <= Pix_326;
    10'd19:  neuron_9_mul_11_p <= Pix_327;
    10'd20:  neuron_9_mul_11_p <= Pix_328;
    10'd21:  neuron_9_mul_11_p <= Pix_329;
    10'd22:  neuron_9_mul_11_p <= Pix_330;
    10'd23:  neuron_9_mul_11_p <= Pix_331;
    10'd24:  neuron_9_mul_11_p <= Pix_332;
    10'd25:  neuron_9_mul_11_p <= Pix_333;
    10'd26:  neuron_9_mul_11_p <= Pix_334;
    10'd27:  neuron_9_mul_11_p <= Pix_335;
    default: neuron_9_mul_11_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_12_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_12_p <= Pix_336;
    10'd1:  neuron_9_mul_12_p <= Pix_337;
    10'd2:  neuron_9_mul_12_p <= Pix_338;
    10'd3:  neuron_9_mul_12_p <= Pix_339;
    10'd4:  neuron_9_mul_12_p <= Pix_340;
    10'd5:  neuron_9_mul_12_p <= Pix_341;
    10'd6:  neuron_9_mul_12_p <= Pix_342;
    10'd7:  neuron_9_mul_12_p <= Pix_343;
    10'd8:  neuron_9_mul_12_p <= Pix_344;
    10'd9:  neuron_9_mul_12_p <= Pix_345;
    10'd10:  neuron_9_mul_12_p <= Pix_346;
    10'd11:  neuron_9_mul_12_p <= Pix_347;
    10'd12:  neuron_9_mul_12_p <= Pix_348;
    10'd13:  neuron_9_mul_12_p <= Pix_349;
    10'd14:  neuron_9_mul_12_p <= Pix_350;
    10'd15:  neuron_9_mul_12_p <= Pix_351;
    10'd16:  neuron_9_mul_12_p <= Pix_352;
    10'd17:  neuron_9_mul_12_p <= Pix_353;
    10'd18:  neuron_9_mul_12_p <= Pix_354;
    10'd19:  neuron_9_mul_12_p <= Pix_355;
    10'd20:  neuron_9_mul_12_p <= Pix_356;
    10'd21:  neuron_9_mul_12_p <= Pix_357;
    10'd22:  neuron_9_mul_12_p <= Pix_358;
    10'd23:  neuron_9_mul_12_p <= Pix_359;
    10'd24:  neuron_9_mul_12_p <= Pix_360;
    10'd25:  neuron_9_mul_12_p <= Pix_361;
    10'd26:  neuron_9_mul_12_p <= Pix_362;
    10'd27:  neuron_9_mul_12_p <= Pix_363;
    default: neuron_9_mul_12_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_13_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_13_p <= Pix_364;
    10'd1:  neuron_9_mul_13_p <= Pix_365;
    10'd2:  neuron_9_mul_13_p <= Pix_366;
    10'd3:  neuron_9_mul_13_p <= Pix_367;
    10'd4:  neuron_9_mul_13_p <= Pix_368;
    10'd5:  neuron_9_mul_13_p <= Pix_369;
    10'd6:  neuron_9_mul_13_p <= Pix_370;
    10'd7:  neuron_9_mul_13_p <= Pix_371;
    10'd8:  neuron_9_mul_13_p <= Pix_372;
    10'd9:  neuron_9_mul_13_p <= Pix_373;
    10'd10:  neuron_9_mul_13_p <= Pix_374;
    10'd11:  neuron_9_mul_13_p <= Pix_375;
    10'd12:  neuron_9_mul_13_p <= Pix_376;
    10'd13:  neuron_9_mul_13_p <= Pix_377;
    10'd14:  neuron_9_mul_13_p <= Pix_378;
    10'd15:  neuron_9_mul_13_p <= Pix_379;
    10'd16:  neuron_9_mul_13_p <= Pix_380;
    10'd17:  neuron_9_mul_13_p <= Pix_381;
    10'd18:  neuron_9_mul_13_p <= Pix_382;
    10'd19:  neuron_9_mul_13_p <= Pix_383;
    10'd20:  neuron_9_mul_13_p <= Pix_384;
    10'd21:  neuron_9_mul_13_p <= Pix_385;
    10'd22:  neuron_9_mul_13_p <= Pix_386;
    10'd23:  neuron_9_mul_13_p <= Pix_387;
    10'd24:  neuron_9_mul_13_p <= Pix_388;
    10'd25:  neuron_9_mul_13_p <= Pix_389;
    10'd26:  neuron_9_mul_13_p <= Pix_390;
    10'd27:  neuron_9_mul_13_p <= Pix_391;
    default: neuron_9_mul_13_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_14_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_14_p <= Pix_392;
    10'd1:  neuron_9_mul_14_p <= Pix_393;
    10'd2:  neuron_9_mul_14_p <= Pix_394;
    10'd3:  neuron_9_mul_14_p <= Pix_395;
    10'd4:  neuron_9_mul_14_p <= Pix_396;
    10'd5:  neuron_9_mul_14_p <= Pix_397;
    10'd6:  neuron_9_mul_14_p <= Pix_398;
    10'd7:  neuron_9_mul_14_p <= Pix_399;
    10'd8:  neuron_9_mul_14_p <= Pix_400;
    10'd9:  neuron_9_mul_14_p <= Pix_401;
    10'd10:  neuron_9_mul_14_p <= Pix_402;
    10'd11:  neuron_9_mul_14_p <= Pix_403;
    10'd12:  neuron_9_mul_14_p <= Pix_404;
    10'd13:  neuron_9_mul_14_p <= Pix_405;
    10'd14:  neuron_9_mul_14_p <= Pix_406;
    10'd15:  neuron_9_mul_14_p <= Pix_407;
    10'd16:  neuron_9_mul_14_p <= Pix_408;
    10'd17:  neuron_9_mul_14_p <= Pix_409;
    10'd18:  neuron_9_mul_14_p <= Pix_410;
    10'd19:  neuron_9_mul_14_p <= Pix_411;
    10'd20:  neuron_9_mul_14_p <= Pix_412;
    10'd21:  neuron_9_mul_14_p <= Pix_413;
    10'd22:  neuron_9_mul_14_p <= Pix_414;
    10'd23:  neuron_9_mul_14_p <= Pix_415;
    10'd24:  neuron_9_mul_14_p <= Pix_416;
    10'd25:  neuron_9_mul_14_p <= Pix_417;
    10'd26:  neuron_9_mul_14_p <= Pix_418;
    10'd27:  neuron_9_mul_14_p <= Pix_419;
    default: neuron_9_mul_14_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_15_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_15_p <= Pix_420;
    10'd1:  neuron_9_mul_15_p <= Pix_421;
    10'd2:  neuron_9_mul_15_p <= Pix_422;
    10'd3:  neuron_9_mul_15_p <= Pix_423;
    10'd4:  neuron_9_mul_15_p <= Pix_424;
    10'd5:  neuron_9_mul_15_p <= Pix_425;
    10'd6:  neuron_9_mul_15_p <= Pix_426;
    10'd7:  neuron_9_mul_15_p <= Pix_427;
    10'd8:  neuron_9_mul_15_p <= Pix_428;
    10'd9:  neuron_9_mul_15_p <= Pix_429;
    10'd10:  neuron_9_mul_15_p <= Pix_430;
    10'd11:  neuron_9_mul_15_p <= Pix_431;
    10'd12:  neuron_9_mul_15_p <= Pix_432;
    10'd13:  neuron_9_mul_15_p <= Pix_433;
    10'd14:  neuron_9_mul_15_p <= Pix_434;
    10'd15:  neuron_9_mul_15_p <= Pix_435;
    10'd16:  neuron_9_mul_15_p <= Pix_436;
    10'd17:  neuron_9_mul_15_p <= Pix_437;
    10'd18:  neuron_9_mul_15_p <= Pix_438;
    10'd19:  neuron_9_mul_15_p <= Pix_439;
    10'd20:  neuron_9_mul_15_p <= Pix_440;
    10'd21:  neuron_9_mul_15_p <= Pix_441;
    10'd22:  neuron_9_mul_15_p <= Pix_442;
    10'd23:  neuron_9_mul_15_p <= Pix_443;
    10'd24:  neuron_9_mul_15_p <= Pix_444;
    10'd25:  neuron_9_mul_15_p <= Pix_445;
    10'd26:  neuron_9_mul_15_p <= Pix_446;
    10'd27:  neuron_9_mul_15_p <= Pix_447;
    default: neuron_9_mul_15_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_16_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_16_p <= Pix_448;
    10'd1:  neuron_9_mul_16_p <= Pix_449;
    10'd2:  neuron_9_mul_16_p <= Pix_450;
    10'd3:  neuron_9_mul_16_p <= Pix_451;
    10'd4:  neuron_9_mul_16_p <= Pix_452;
    10'd5:  neuron_9_mul_16_p <= Pix_453;
    10'd6:  neuron_9_mul_16_p <= Pix_454;
    10'd7:  neuron_9_mul_16_p <= Pix_455;
    10'd8:  neuron_9_mul_16_p <= Pix_456;
    10'd9:  neuron_9_mul_16_p <= Pix_457;
    10'd10:  neuron_9_mul_16_p <= Pix_458;
    10'd11:  neuron_9_mul_16_p <= Pix_459;
    10'd12:  neuron_9_mul_16_p <= Pix_460;
    10'd13:  neuron_9_mul_16_p <= Pix_461;
    10'd14:  neuron_9_mul_16_p <= Pix_462;
    10'd15:  neuron_9_mul_16_p <= Pix_463;
    10'd16:  neuron_9_mul_16_p <= Pix_464;
    10'd17:  neuron_9_mul_16_p <= Pix_465;
    10'd18:  neuron_9_mul_16_p <= Pix_466;
    10'd19:  neuron_9_mul_16_p <= Pix_467;
    10'd20:  neuron_9_mul_16_p <= Pix_468;
    10'd21:  neuron_9_mul_16_p <= Pix_469;
    10'd22:  neuron_9_mul_16_p <= Pix_470;
    10'd23:  neuron_9_mul_16_p <= Pix_471;
    10'd24:  neuron_9_mul_16_p <= Pix_472;
    10'd25:  neuron_9_mul_16_p <= Pix_473;
    10'd26:  neuron_9_mul_16_p <= Pix_474;
    10'd27:  neuron_9_mul_16_p <= Pix_475;
    default: neuron_9_mul_16_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_17_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_17_p <= Pix_476;
    10'd1:  neuron_9_mul_17_p <= Pix_477;
    10'd2:  neuron_9_mul_17_p <= Pix_478;
    10'd3:  neuron_9_mul_17_p <= Pix_479;
    10'd4:  neuron_9_mul_17_p <= Pix_480;
    10'd5:  neuron_9_mul_17_p <= Pix_481;
    10'd6:  neuron_9_mul_17_p <= Pix_482;
    10'd7:  neuron_9_mul_17_p <= Pix_483;
    10'd8:  neuron_9_mul_17_p <= Pix_484;
    10'd9:  neuron_9_mul_17_p <= Pix_485;
    10'd10:  neuron_9_mul_17_p <= Pix_486;
    10'd11:  neuron_9_mul_17_p <= Pix_487;
    10'd12:  neuron_9_mul_17_p <= Pix_488;
    10'd13:  neuron_9_mul_17_p <= Pix_489;
    10'd14:  neuron_9_mul_17_p <= Pix_490;
    10'd15:  neuron_9_mul_17_p <= Pix_491;
    10'd16:  neuron_9_mul_17_p <= Pix_492;
    10'd17:  neuron_9_mul_17_p <= Pix_493;
    10'd18:  neuron_9_mul_17_p <= Pix_494;
    10'd19:  neuron_9_mul_17_p <= Pix_495;
    10'd20:  neuron_9_mul_17_p <= Pix_496;
    10'd21:  neuron_9_mul_17_p <= Pix_497;
    10'd22:  neuron_9_mul_17_p <= Pix_498;
    10'd23:  neuron_9_mul_17_p <= Pix_499;
    10'd24:  neuron_9_mul_17_p <= Pix_500;
    10'd25:  neuron_9_mul_17_p <= Pix_501;
    10'd26:  neuron_9_mul_17_p <= Pix_502;
    10'd27:  neuron_9_mul_17_p <= Pix_503;
    default: neuron_9_mul_17_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_18_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_18_p <= Pix_504;
    10'd1:  neuron_9_mul_18_p <= Pix_505;
    10'd2:  neuron_9_mul_18_p <= Pix_506;
    10'd3:  neuron_9_mul_18_p <= Pix_507;
    10'd4:  neuron_9_mul_18_p <= Pix_508;
    10'd5:  neuron_9_mul_18_p <= Pix_509;
    10'd6:  neuron_9_mul_18_p <= Pix_510;
    10'd7:  neuron_9_mul_18_p <= Pix_511;
    10'd8:  neuron_9_mul_18_p <= Pix_512;
    10'd9:  neuron_9_mul_18_p <= Pix_513;
    10'd10:  neuron_9_mul_18_p <= Pix_514;
    10'd11:  neuron_9_mul_18_p <= Pix_515;
    10'd12:  neuron_9_mul_18_p <= Pix_516;
    10'd13:  neuron_9_mul_18_p <= Pix_517;
    10'd14:  neuron_9_mul_18_p <= Pix_518;
    10'd15:  neuron_9_mul_18_p <= Pix_519;
    10'd16:  neuron_9_mul_18_p <= Pix_520;
    10'd17:  neuron_9_mul_18_p <= Pix_521;
    10'd18:  neuron_9_mul_18_p <= Pix_522;
    10'd19:  neuron_9_mul_18_p <= Pix_523;
    10'd20:  neuron_9_mul_18_p <= Pix_524;
    10'd21:  neuron_9_mul_18_p <= Pix_525;
    10'd22:  neuron_9_mul_18_p <= Pix_526;
    10'd23:  neuron_9_mul_18_p <= Pix_527;
    10'd24:  neuron_9_mul_18_p <= Pix_528;
    10'd25:  neuron_9_mul_18_p <= Pix_529;
    10'd26:  neuron_9_mul_18_p <= Pix_530;
    10'd27:  neuron_9_mul_18_p <= Pix_531;
    default: neuron_9_mul_18_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_19_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_19_p <= Pix_532;
    10'd1:  neuron_9_mul_19_p <= Pix_533;
    10'd2:  neuron_9_mul_19_p <= Pix_534;
    10'd3:  neuron_9_mul_19_p <= Pix_535;
    10'd4:  neuron_9_mul_19_p <= Pix_536;
    10'd5:  neuron_9_mul_19_p <= Pix_537;
    10'd6:  neuron_9_mul_19_p <= Pix_538;
    10'd7:  neuron_9_mul_19_p <= Pix_539;
    10'd8:  neuron_9_mul_19_p <= Pix_540;
    10'd9:  neuron_9_mul_19_p <= Pix_541;
    10'd10:  neuron_9_mul_19_p <= Pix_542;
    10'd11:  neuron_9_mul_19_p <= Pix_543;
    10'd12:  neuron_9_mul_19_p <= Pix_544;
    10'd13:  neuron_9_mul_19_p <= Pix_545;
    10'd14:  neuron_9_mul_19_p <= Pix_546;
    10'd15:  neuron_9_mul_19_p <= Pix_547;
    10'd16:  neuron_9_mul_19_p <= Pix_548;
    10'd17:  neuron_9_mul_19_p <= Pix_549;
    10'd18:  neuron_9_mul_19_p <= Pix_550;
    10'd19:  neuron_9_mul_19_p <= Pix_551;
    10'd20:  neuron_9_mul_19_p <= Pix_552;
    10'd21:  neuron_9_mul_19_p <= Pix_553;
    10'd22:  neuron_9_mul_19_p <= Pix_554;
    10'd23:  neuron_9_mul_19_p <= Pix_555;
    10'd24:  neuron_9_mul_19_p <= Pix_556;
    10'd25:  neuron_9_mul_19_p <= Pix_557;
    10'd26:  neuron_9_mul_19_p <= Pix_558;
    10'd27:  neuron_9_mul_19_p <= Pix_559;
    default: neuron_9_mul_19_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_20_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_20_p <= Pix_560;
    10'd1:  neuron_9_mul_20_p <= Pix_561;
    10'd2:  neuron_9_mul_20_p <= Pix_562;
    10'd3:  neuron_9_mul_20_p <= Pix_563;
    10'd4:  neuron_9_mul_20_p <= Pix_564;
    10'd5:  neuron_9_mul_20_p <= Pix_565;
    10'd6:  neuron_9_mul_20_p <= Pix_566;
    10'd7:  neuron_9_mul_20_p <= Pix_567;
    10'd8:  neuron_9_mul_20_p <= Pix_568;
    10'd9:  neuron_9_mul_20_p <= Pix_569;
    10'd10:  neuron_9_mul_20_p <= Pix_570;
    10'd11:  neuron_9_mul_20_p <= Pix_571;
    10'd12:  neuron_9_mul_20_p <= Pix_572;
    10'd13:  neuron_9_mul_20_p <= Pix_573;
    10'd14:  neuron_9_mul_20_p <= Pix_574;
    10'd15:  neuron_9_mul_20_p <= Pix_575;
    10'd16:  neuron_9_mul_20_p <= Pix_576;
    10'd17:  neuron_9_mul_20_p <= Pix_577;
    10'd18:  neuron_9_mul_20_p <= Pix_578;
    10'd19:  neuron_9_mul_20_p <= Pix_579;
    10'd20:  neuron_9_mul_20_p <= Pix_580;
    10'd21:  neuron_9_mul_20_p <= Pix_581;
    10'd22:  neuron_9_mul_20_p <= Pix_582;
    10'd23:  neuron_9_mul_20_p <= Pix_583;
    10'd24:  neuron_9_mul_20_p <= Pix_584;
    10'd25:  neuron_9_mul_20_p <= Pix_585;
    10'd26:  neuron_9_mul_20_p <= Pix_586;
    10'd27:  neuron_9_mul_20_p <= Pix_587;
    default: neuron_9_mul_20_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_21_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_21_p <= Pix_588;
    10'd1:  neuron_9_mul_21_p <= Pix_589;
    10'd2:  neuron_9_mul_21_p <= Pix_590;
    10'd3:  neuron_9_mul_21_p <= Pix_591;
    10'd4:  neuron_9_mul_21_p <= Pix_592;
    10'd5:  neuron_9_mul_21_p <= Pix_593;
    10'd6:  neuron_9_mul_21_p <= Pix_594;
    10'd7:  neuron_9_mul_21_p <= Pix_595;
    10'd8:  neuron_9_mul_21_p <= Pix_596;
    10'd9:  neuron_9_mul_21_p <= Pix_597;
    10'd10:  neuron_9_mul_21_p <= Pix_598;
    10'd11:  neuron_9_mul_21_p <= Pix_599;
    10'd12:  neuron_9_mul_21_p <= Pix_600;
    10'd13:  neuron_9_mul_21_p <= Pix_601;
    10'd14:  neuron_9_mul_21_p <= Pix_602;
    10'd15:  neuron_9_mul_21_p <= Pix_603;
    10'd16:  neuron_9_mul_21_p <= Pix_604;
    10'd17:  neuron_9_mul_21_p <= Pix_605;
    10'd18:  neuron_9_mul_21_p <= Pix_606;
    10'd19:  neuron_9_mul_21_p <= Pix_607;
    10'd20:  neuron_9_mul_21_p <= Pix_608;
    10'd21:  neuron_9_mul_21_p <= Pix_609;
    10'd22:  neuron_9_mul_21_p <= Pix_610;
    10'd23:  neuron_9_mul_21_p <= Pix_611;
    10'd24:  neuron_9_mul_21_p <= Pix_612;
    10'd25:  neuron_9_mul_21_p <= Pix_613;
    10'd26:  neuron_9_mul_21_p <= Pix_614;
    10'd27:  neuron_9_mul_21_p <= Pix_615;
    default: neuron_9_mul_21_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_22_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_22_p <= Pix_616;
    10'd1:  neuron_9_mul_22_p <= Pix_617;
    10'd2:  neuron_9_mul_22_p <= Pix_618;
    10'd3:  neuron_9_mul_22_p <= Pix_619;
    10'd4:  neuron_9_mul_22_p <= Pix_620;
    10'd5:  neuron_9_mul_22_p <= Pix_621;
    10'd6:  neuron_9_mul_22_p <= Pix_622;
    10'd7:  neuron_9_mul_22_p <= Pix_623;
    10'd8:  neuron_9_mul_22_p <= Pix_624;
    10'd9:  neuron_9_mul_22_p <= Pix_625;
    10'd10:  neuron_9_mul_22_p <= Pix_626;
    10'd11:  neuron_9_mul_22_p <= Pix_627;
    10'd12:  neuron_9_mul_22_p <= Pix_628;
    10'd13:  neuron_9_mul_22_p <= Pix_629;
    10'd14:  neuron_9_mul_22_p <= Pix_630;
    10'd15:  neuron_9_mul_22_p <= Pix_631;
    10'd16:  neuron_9_mul_22_p <= Pix_632;
    10'd17:  neuron_9_mul_22_p <= Pix_633;
    10'd18:  neuron_9_mul_22_p <= Pix_634;
    10'd19:  neuron_9_mul_22_p <= Pix_635;
    10'd20:  neuron_9_mul_22_p <= Pix_636;
    10'd21:  neuron_9_mul_22_p <= Pix_637;
    10'd22:  neuron_9_mul_22_p <= Pix_638;
    10'd23:  neuron_9_mul_22_p <= Pix_639;
    10'd24:  neuron_9_mul_22_p <= Pix_640;
    10'd25:  neuron_9_mul_22_p <= Pix_641;
    10'd26:  neuron_9_mul_22_p <= Pix_642;
    10'd27:  neuron_9_mul_22_p <= Pix_643;
    default: neuron_9_mul_22_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_23_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_23_p <= Pix_644;
    10'd1:  neuron_9_mul_23_p <= Pix_645;
    10'd2:  neuron_9_mul_23_p <= Pix_646;
    10'd3:  neuron_9_mul_23_p <= Pix_647;
    10'd4:  neuron_9_mul_23_p <= Pix_648;
    10'd5:  neuron_9_mul_23_p <= Pix_649;
    10'd6:  neuron_9_mul_23_p <= Pix_650;
    10'd7:  neuron_9_mul_23_p <= Pix_651;
    10'd8:  neuron_9_mul_23_p <= Pix_652;
    10'd9:  neuron_9_mul_23_p <= Pix_653;
    10'd10:  neuron_9_mul_23_p <= Pix_654;
    10'd11:  neuron_9_mul_23_p <= Pix_655;
    10'd12:  neuron_9_mul_23_p <= Pix_656;
    10'd13:  neuron_9_mul_23_p <= Pix_657;
    10'd14:  neuron_9_mul_23_p <= Pix_658;
    10'd15:  neuron_9_mul_23_p <= Pix_659;
    10'd16:  neuron_9_mul_23_p <= Pix_660;
    10'd17:  neuron_9_mul_23_p <= Pix_661;
    10'd18:  neuron_9_mul_23_p <= Pix_662;
    10'd19:  neuron_9_mul_23_p <= Pix_663;
    10'd20:  neuron_9_mul_23_p <= Pix_664;
    10'd21:  neuron_9_mul_23_p <= Pix_665;
    10'd22:  neuron_9_mul_23_p <= Pix_666;
    10'd23:  neuron_9_mul_23_p <= Pix_667;
    10'd24:  neuron_9_mul_23_p <= Pix_668;
    10'd25:  neuron_9_mul_23_p <= Pix_669;
    10'd26:  neuron_9_mul_23_p <= Pix_670;
    10'd27:  neuron_9_mul_23_p <= Pix_671;
    default: neuron_9_mul_23_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_24_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_24_p <= Pix_672;
    10'd1:  neuron_9_mul_24_p <= Pix_673;
    10'd2:  neuron_9_mul_24_p <= Pix_674;
    10'd3:  neuron_9_mul_24_p <= Pix_675;
    10'd4:  neuron_9_mul_24_p <= Pix_676;
    10'd5:  neuron_9_mul_24_p <= Pix_677;
    10'd6:  neuron_9_mul_24_p <= Pix_678;
    10'd7:  neuron_9_mul_24_p <= Pix_679;
    10'd8:  neuron_9_mul_24_p <= Pix_680;
    10'd9:  neuron_9_mul_24_p <= Pix_681;
    10'd10:  neuron_9_mul_24_p <= Pix_682;
    10'd11:  neuron_9_mul_24_p <= Pix_683;
    10'd12:  neuron_9_mul_24_p <= Pix_684;
    10'd13:  neuron_9_mul_24_p <= Pix_685;
    10'd14:  neuron_9_mul_24_p <= Pix_686;
    10'd15:  neuron_9_mul_24_p <= Pix_687;
    10'd16:  neuron_9_mul_24_p <= Pix_688;
    10'd17:  neuron_9_mul_24_p <= Pix_689;
    10'd18:  neuron_9_mul_24_p <= Pix_690;
    10'd19:  neuron_9_mul_24_p <= Pix_691;
    10'd20:  neuron_9_mul_24_p <= Pix_692;
    10'd21:  neuron_9_mul_24_p <= Pix_693;
    10'd22:  neuron_9_mul_24_p <= Pix_694;
    10'd23:  neuron_9_mul_24_p <= Pix_695;
    10'd24:  neuron_9_mul_24_p <= Pix_696;
    10'd25:  neuron_9_mul_24_p <= Pix_697;
    10'd26:  neuron_9_mul_24_p <= Pix_698;
    10'd27:  neuron_9_mul_24_p <= Pix_699;
    default: neuron_9_mul_24_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_25_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_25_p <= Pix_700;
    10'd1:  neuron_9_mul_25_p <= Pix_701;
    10'd2:  neuron_9_mul_25_p <= Pix_702;
    10'd3:  neuron_9_mul_25_p <= Pix_703;
    10'd4:  neuron_9_mul_25_p <= Pix_704;
    10'd5:  neuron_9_mul_25_p <= Pix_705;
    10'd6:  neuron_9_mul_25_p <= Pix_706;
    10'd7:  neuron_9_mul_25_p <= Pix_707;
    10'd8:  neuron_9_mul_25_p <= Pix_708;
    10'd9:  neuron_9_mul_25_p <= Pix_709;
    10'd10:  neuron_9_mul_25_p <= Pix_710;
    10'd11:  neuron_9_mul_25_p <= Pix_711;
    10'd12:  neuron_9_mul_25_p <= Pix_712;
    10'd13:  neuron_9_mul_25_p <= Pix_713;
    10'd14:  neuron_9_mul_25_p <= Pix_714;
    10'd15:  neuron_9_mul_25_p <= Pix_715;
    10'd16:  neuron_9_mul_25_p <= Pix_716;
    10'd17:  neuron_9_mul_25_p <= Pix_717;
    10'd18:  neuron_9_mul_25_p <= Pix_718;
    10'd19:  neuron_9_mul_25_p <= Pix_719;
    10'd20:  neuron_9_mul_25_p <= Pix_720;
    10'd21:  neuron_9_mul_25_p <= Pix_721;
    10'd22:  neuron_9_mul_25_p <= Pix_722;
    10'd23:  neuron_9_mul_25_p <= Pix_723;
    10'd24:  neuron_9_mul_25_p <= Pix_724;
    10'd25:  neuron_9_mul_25_p <= Pix_725;
    10'd26:  neuron_9_mul_25_p <= Pix_726;
    10'd27:  neuron_9_mul_25_p <= Pix_727;
    default: neuron_9_mul_25_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_26_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_26_p <= Pix_728;
    10'd1:  neuron_9_mul_26_p <= Pix_729;
    10'd2:  neuron_9_mul_26_p <= Pix_730;
    10'd3:  neuron_9_mul_26_p <= Pix_731;
    10'd4:  neuron_9_mul_26_p <= Pix_732;
    10'd5:  neuron_9_mul_26_p <= Pix_733;
    10'd6:  neuron_9_mul_26_p <= Pix_734;
    10'd7:  neuron_9_mul_26_p <= Pix_735;
    10'd8:  neuron_9_mul_26_p <= Pix_736;
    10'd9:  neuron_9_mul_26_p <= Pix_737;
    10'd10:  neuron_9_mul_26_p <= Pix_738;
    10'd11:  neuron_9_mul_26_p <= Pix_739;
    10'd12:  neuron_9_mul_26_p <= Pix_740;
    10'd13:  neuron_9_mul_26_p <= Pix_741;
    10'd14:  neuron_9_mul_26_p <= Pix_742;
    10'd15:  neuron_9_mul_26_p <= Pix_743;
    10'd16:  neuron_9_mul_26_p <= Pix_744;
    10'd17:  neuron_9_mul_26_p <= Pix_745;
    10'd18:  neuron_9_mul_26_p <= Pix_746;
    10'd19:  neuron_9_mul_26_p <= Pix_747;
    10'd20:  neuron_9_mul_26_p <= Pix_748;
    10'd21:  neuron_9_mul_26_p <= Pix_749;
    10'd22:  neuron_9_mul_26_p <= Pix_750;
    10'd23:  neuron_9_mul_26_p <= Pix_751;
    10'd24:  neuron_9_mul_26_p <= Pix_752;
    10'd25:  neuron_9_mul_26_p <= Pix_753;
    10'd26:  neuron_9_mul_26_p <= Pix_754;
    10'd27:  neuron_9_mul_26_p <= Pix_755;
    default: neuron_9_mul_26_p <= 0;
  endcase
  end
end

always @(posedge clk) begin
  if(GlobalReset)
    neuron_9_mul_27_p <= 0;
  else begin
  case(N):
    10'd0:  neuron_9_mul_27_p <= Pix_756;
    10'd1:  neuron_9_mul_27_p <= Pix_757;
    10'd2:  neuron_9_mul_27_p <= Pix_758;
    10'd3:  neuron_9_mul_27_p <= Pix_759;
    10'd4:  neuron_9_mul_27_p <= Pix_760;
    10'd5:  neuron_9_mul_27_p <= Pix_761;
    10'd6:  neuron_9_mul_27_p <= Pix_762;
    10'd7:  neuron_9_mul_27_p <= Pix_763;
    10'd8:  neuron_9_mul_27_p <= Pix_764;
    10'd9:  neuron_9_mul_27_p <= Pix_765;
    10'd10:  neuron_9_mul_27_p <= Pix_766;
    10'd11:  neuron_9_mul_27_p <= Pix_767;
    10'd12:  neuron_9_mul_27_p <= Pix_768;
    10'd13:  neuron_9_mul_27_p <= Pix_769;
    10'd14:  neuron_9_mul_27_p <= Pix_770;
    10'd15:  neuron_9_mul_27_p <= Pix_771;
    10'd16:  neuron_9_mul_27_p <= Pix_772;
    10'd17:  neuron_9_mul_27_p <= Pix_773;
    10'd18:  neuron_9_mul_27_p <= Pix_774;
    10'd19:  neuron_9_mul_27_p <= Pix_775;
    10'd20:  neuron_9_mul_27_p <= Pix_776;
    10'd21:  neuron_9_mul_27_p <= Pix_777;
    10'd22:  neuron_9_mul_27_p <= Pix_778;
    10'd23:  neuron_9_mul_27_p <= Pix_779;
    10'd24:  neuron_9_mul_27_p <= Pix_780;
    10'd25:  neuron_9_mul_27_p <= Pix_781;
    10'd26:  neuron_9_mul_27_p <= Pix_782;
    10'd27:  neuron_9_mul_27_p <= Pix_783;
    default: neuron_9_mul_27_p <= 0;
  endcase
  end
end

endmodule
