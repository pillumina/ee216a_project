// Weight: 最高位不是符号位,小数点后18位,即Weight绝对值小于1. 0~0.25
// Pixel: 10位,为什么要10位???! 8位都够了
// V1.0
// For multipliers, its 28*28(bits)*10, 280 multipliers in total
// For adders, its 28*10, 280 in total
// In total, there are 10 neurons and each neuron has 28 multipliers and 28 adders

module Image_Classifier (
 input clk,
 input GlobalReset,   // Apply synchronous active-high reset to all blocks
 input Input_Valid,
 input [18:0] Wgt_0_0, // sfix19_En18
  input [18:0] Wgt_0_1, // sfix19_En18
  input [18:0] Wgt_0_2, // sfix19_En18
  input [18:0] Wgt_0_3, // sfix19_En18
  input [18:0] Wgt_0_4, // sfix19_En18
  input [18:0] Wgt_0_5, // sfix19_En18
  input [18:0] Wgt_0_6, // sfix19_En18
  input [18:0] Wgt_0_7, // sfix19_En18
  input [18:0] Wgt_0_8, // sfix19_En18
  input [18:0] Wgt_0_9, // sfix19_En18
  input [18:0] Wgt_0_10, // sfix19_En18
  input [18:0] Wgt_0_11, // sfix19_En18
  input [18:0] Wgt_0_12, // sfix19_En18
  input [18:0] Wgt_0_13, // sfix19_En18
  input [18:0] Wgt_0_14, // sfix19_En18
  input [18:0] Wgt_0_15, // sfix19_En18
  input [18:0] Wgt_0_16, // sfix19_En18
  input [18:0] Wgt_0_17, // sfix19_En18
  input [18:0] Wgt_0_18, // sfix19_En18
  input [18:0] Wgt_0_19, // sfix19_En18
  input [18:0] Wgt_0_20, // sfix19_En18
  input [18:0] Wgt_0_21, // sfix19_En18
  input [18:0] Wgt_0_22, // sfix19_En18
  input [18:0] Wgt_0_23, // sfix19_En18
  input [18:0] Wgt_0_24, // sfix19_En18
  input [18:0] Wgt_0_25, // sfix19_En18
  input [18:0] Wgt_0_26, // sfix19_En18
  input [18:0] Wgt_0_27, // sfix19_En18
  input [18:0] Wgt_0_28, // sfix19_En18
  input [18:0] Wgt_0_29, // sfix19_En18
  input [18:0] Wgt_0_30, // sfix19_En18
  input [18:0] Wgt_0_31, // sfix19_En18
  input [18:0] Wgt_0_32, // sfix19_En18
  input [18:0] Wgt_0_33, // sfix19_En18
  input [18:0] Wgt_0_34, // sfix19_En18
  input [18:0] Wgt_0_35, // sfix19_En18
  input [18:0] Wgt_0_36, // sfix19_En18
  input [18:0] Wgt_0_37, // sfix19_En18
  input [18:0] Wgt_0_38, // sfix19_En18
  input [18:0] Wgt_0_39, // sfix19_En18
  input [18:0] Wgt_0_40, // sfix19_En18
  input [18:0] Wgt_0_41, // sfix19_En18
  input [18:0] Wgt_0_42, // sfix19_En18
  input [18:0] Wgt_0_43, // sfix19_En18
  input [18:0] Wgt_0_44, // sfix19_En18
  input [18:0] Wgt_0_45, // sfix19_En18
  input [18:0] Wgt_0_46, // sfix19_En18
  input [18:0] Wgt_0_47, // sfix19_En18
  input [18:0] Wgt_0_48, // sfix19_En18
  input [18:0] Wgt_0_49, // sfix19_En18
  input [18:0] Wgt_0_50, // sfix19_En18
  input [18:0] Wgt_0_51, // sfix19_En18
  input [18:0] Wgt_0_52, // sfix19_En18
  input [18:0] Wgt_0_53, // sfix19_En18
  input [18:0] Wgt_0_54, // sfix19_En18
  input [18:0] Wgt_0_55, // sfix19_En18
  input [18:0] Wgt_0_56, // sfix19_En18
  input [18:0] Wgt_0_57, // sfix19_En18
  input [18:0] Wgt_0_58, // sfix19_En18
  input [18:0] Wgt_0_59, // sfix19_En18
  input [18:0] Wgt_0_60, // sfix19_En18
  input [18:0] Wgt_0_61, // sfix19_En18
  input [18:0] Wgt_0_62, // sfix19_En18
  input [18:0] Wgt_0_63, // sfix19_En18
  input [18:0] Wgt_0_64, // sfix19_En18
  input [18:0] Wgt_0_65, // sfix19_En18
  input [18:0] Wgt_0_66, // sfix19_En18
  input [18:0] Wgt_0_67, // sfix19_En18
  input [18:0] Wgt_0_68, // sfix19_En18
  input [18:0] Wgt_0_69, // sfix19_En18
  input [18:0] Wgt_0_70, // sfix19_En18
  input [18:0] Wgt_0_71, // sfix19_En18
  input [18:0] Wgt_0_72, // sfix19_En18
  input [18:0] Wgt_0_73, // sfix19_En18
  input [18:0] Wgt_0_74, // sfix19_En18
  input [18:0] Wgt_0_75, // sfix19_En18
  input [18:0] Wgt_0_76, // sfix19_En18
  input [18:0] Wgt_0_77, // sfix19_En18
  input [18:0] Wgt_0_78, // sfix19_En18
  input [18:0] Wgt_0_79, // sfix19_En18
  input [18:0] Wgt_0_80, // sfix19_En18
  input [18:0] Wgt_0_81, // sfix19_En18
  input [18:0] Wgt_0_82, // sfix19_En18
  input [18:0] Wgt_0_83, // sfix19_En18
  input [18:0] Wgt_0_84, // sfix19_En18
  input [18:0] Wgt_0_85, // sfix19_En18
  input [18:0] Wgt_0_86, // sfix19_En18
  input [18:0] Wgt_0_87, // sfix19_En18
  input [18:0] Wgt_0_88, // sfix19_En18
  input [18:0] Wgt_0_89, // sfix19_En18
  input [18:0] Wgt_0_90, // sfix19_En18
  input [18:0] Wgt_0_91, // sfix19_En18
  input [18:0] Wgt_0_92, // sfix19_En18
  input [18:0] Wgt_0_93, // sfix19_En18
  input [18:0] Wgt_0_94, // sfix19_En18
  input [18:0] Wgt_0_95, // sfix19_En18
  input [18:0] Wgt_0_96, // sfix19_En18
  input [18:0] Wgt_0_97, // sfix19_En18
  input [18:0] Wgt_0_98, // sfix19_En18
  input [18:0] Wgt_0_99, // sfix19_En18
  input [18:0] Wgt_0_100, // sfix19_En18
  input [18:0] Wgt_0_101, // sfix19_En18
  input [18:0] Wgt_0_102, // sfix19_En18
  input [18:0] Wgt_0_103, // sfix19_En18
  input [18:0] Wgt_0_104, // sfix19_En18
  input [18:0] Wgt_0_105, // sfix19_En18
  input [18:0] Wgt_0_106, // sfix19_En18
  input [18:0] Wgt_0_107, // sfix19_En18
  input [18:0] Wgt_0_108, // sfix19_En18
  input [18:0] Wgt_0_109, // sfix19_En18
  input [18:0] Wgt_0_110, // sfix19_En18
  input [18:0] Wgt_0_111, // sfix19_En18
  input [18:0] Wgt_0_112, // sfix19_En18
  input [18:0] Wgt_0_113, // sfix19_En18
  input [18:0] Wgt_0_114, // sfix19_En18
  input [18:0] Wgt_0_115, // sfix19_En18
  input [18:0] Wgt_0_116, // sfix19_En18
  input [18:0] Wgt_0_117, // sfix19_En18
  input [18:0] Wgt_0_118, // sfix19_En18
  input [18:0] Wgt_0_119, // sfix19_En18
  input [18:0] Wgt_0_120, // sfix19_En18
  input [18:0] Wgt_0_121, // sfix19_En18
  input [18:0] Wgt_0_122, // sfix19_En18
  input [18:0] Wgt_0_123, // sfix19_En18
  input [18:0] Wgt_0_124, // sfix19_En18
  input [18:0] Wgt_0_125, // sfix19_En18
  input [18:0] Wgt_0_126, // sfix19_En18
  input [18:0] Wgt_0_127, // sfix19_En18
  input [18:0] Wgt_0_128, // sfix19_En18
  input [18:0] Wgt_0_129, // sfix19_En18
  input [18:0] Wgt_0_130, // sfix19_En18
  input [18:0] Wgt_0_131, // sfix19_En18
  input [18:0] Wgt_0_132, // sfix19_En18
  input [18:0] Wgt_0_133, // sfix19_En18
  input [18:0] Wgt_0_134, // sfix19_En18
  input [18:0] Wgt_0_135, // sfix19_En18
  input [18:0] Wgt_0_136, // sfix19_En18
  input [18:0] Wgt_0_137, // sfix19_En18
  input [18:0] Wgt_0_138, // sfix19_En18
  input [18:0] Wgt_0_139, // sfix19_En18
  input [18:0] Wgt_0_140, // sfix19_En18
  input [18:0] Wgt_0_141, // sfix19_En18
  input [18:0] Wgt_0_142, // sfix19_En18
  input [18:0] Wgt_0_143, // sfix19_En18
  input [18:0] Wgt_0_144, // sfix19_En18
  input [18:0] Wgt_0_145, // sfix19_En18
  input [18:0] Wgt_0_146, // sfix19_En18
  input [18:0] Wgt_0_147, // sfix19_En18
  input [18:0] Wgt_0_148, // sfix19_En18
  input [18:0] Wgt_0_149, // sfix19_En18
  input [18:0] Wgt_0_150, // sfix19_En18
  input [18:0] Wgt_0_151, // sfix19_En18
  input [18:0] Wgt_0_152, // sfix19_En18
  input [18:0] Wgt_0_153, // sfix19_En18
  input [18:0] Wgt_0_154, // sfix19_En18
  input [18:0] Wgt_0_155, // sfix19_En18
  input [18:0] Wgt_0_156, // sfix19_En18
  input [18:0] Wgt_0_157, // sfix19_En18
  input [18:0] Wgt_0_158, // sfix19_En18
  input [18:0] Wgt_0_159, // sfix19_En18
  input [18:0] Wgt_0_160, // sfix19_En18
  input [18:0] Wgt_0_161, // sfix19_En18
  input [18:0] Wgt_0_162, // sfix19_En18
  input [18:0] Wgt_0_163, // sfix19_En18
  input [18:0] Wgt_0_164, // sfix19_En18
  input [18:0] Wgt_0_165, // sfix19_En18
  input [18:0] Wgt_0_166, // sfix19_En18
  input [18:0] Wgt_0_167, // sfix19_En18
  input [18:0] Wgt_0_168, // sfix19_En18
  input [18:0] Wgt_0_169, // sfix19_En18
  input [18:0] Wgt_0_170, // sfix19_En18
  input [18:0] Wgt_0_171, // sfix19_En18
  input [18:0] Wgt_0_172, // sfix19_En18
  input [18:0] Wgt_0_173, // sfix19_En18
  input [18:0] Wgt_0_174, // sfix19_En18
  input [18:0] Wgt_0_175, // sfix19_En18
  input [18:0] Wgt_0_176, // sfix19_En18
  input [18:0] Wgt_0_177, // sfix19_En18
  input [18:0] Wgt_0_178, // sfix19_En18
  input [18:0] Wgt_0_179, // sfix19_En18
  input [18:0] Wgt_0_180, // sfix19_En18
  input [18:0] Wgt_0_181, // sfix19_En18
  input [18:0] Wgt_0_182, // sfix19_En18
  input [18:0] Wgt_0_183, // sfix19_En18
  input [18:0] Wgt_0_184, // sfix19_En18
  input [18:0] Wgt_0_185, // sfix19_En18
  input [18:0] Wgt_0_186, // sfix19_En18
  input [18:0] Wgt_0_187, // sfix19_En18
  input [18:0] Wgt_0_188, // sfix19_En18
  input [18:0] Wgt_0_189, // sfix19_En18
  input [18:0] Wgt_0_190, // sfix19_En18
  input [18:0] Wgt_0_191, // sfix19_En18
  input [18:0] Wgt_0_192, // sfix19_En18
  input [18:0] Wgt_0_193, // sfix19_En18
  input [18:0] Wgt_0_194, // sfix19_En18
  input [18:0] Wgt_0_195, // sfix19_En18
  input [18:0] Wgt_0_196, // sfix19_En18
  input [18:0] Wgt_0_197, // sfix19_En18
  input [18:0] Wgt_0_198, // sfix19_En18
  input [18:0] Wgt_0_199, // sfix19_En18
  input [18:0] Wgt_0_200, // sfix19_En18
  input [18:0] Wgt_0_201, // sfix19_En18
  input [18:0] Wgt_0_202, // sfix19_En18
  input [18:0] Wgt_0_203, // sfix19_En18
  input [18:0] Wgt_0_204, // sfix19_En18
  input [18:0] Wgt_0_205, // sfix19_En18
  input [18:0] Wgt_0_206, // sfix19_En18
  input [18:0] Wgt_0_207, // sfix19_En18
  input [18:0] Wgt_0_208, // sfix19_En18
  input [18:0] Wgt_0_209, // sfix19_En18
  input [18:0] Wgt_0_210, // sfix19_En18
  input [18:0] Wgt_0_211, // sfix19_En18
  input [18:0] Wgt_0_212, // sfix19_En18
  input [18:0] Wgt_0_213, // sfix19_En18
  input [18:0] Wgt_0_214, // sfix19_En18
  input [18:0] Wgt_0_215, // sfix19_En18
  input [18:0] Wgt_0_216, // sfix19_En18
  input [18:0] Wgt_0_217, // sfix19_En18
  input [18:0] Wgt_0_218, // sfix19_En18
  input [18:0] Wgt_0_219, // sfix19_En18
  input [18:0] Wgt_0_220, // sfix19_En18
  input [18:0] Wgt_0_221, // sfix19_En18
  input [18:0] Wgt_0_222, // sfix19_En18
  input [18:0] Wgt_0_223, // sfix19_En18
  input [18:0] Wgt_0_224, // sfix19_En18
  input [18:0] Wgt_0_225, // sfix19_En18
  input [18:0] Wgt_0_226, // sfix19_En18
  input [18:0] Wgt_0_227, // sfix19_En18
  input [18:0] Wgt_0_228, // sfix19_En18
  input [18:0] Wgt_0_229, // sfix19_En18
  input [18:0] Wgt_0_230, // sfix19_En18
  input [18:0] Wgt_0_231, // sfix19_En18
  input [18:0] Wgt_0_232, // sfix19_En18
  input [18:0] Wgt_0_233, // sfix19_En18
  input [18:0] Wgt_0_234, // sfix19_En18
  input [18:0] Wgt_0_235, // sfix19_En18
  input [18:0] Wgt_0_236, // sfix19_En18
  input [18:0] Wgt_0_237, // sfix19_En18
  input [18:0] Wgt_0_238, // sfix19_En18
  input [18:0] Wgt_0_239, // sfix19_En18
  input [18:0] Wgt_0_240, // sfix19_En18
  input [18:0] Wgt_0_241, // sfix19_En18
  input [18:0] Wgt_0_242, // sfix19_En18
  input [18:0] Wgt_0_243, // sfix19_En18
  input [18:0] Wgt_0_244, // sfix19_En18
  input [18:0] Wgt_0_245, // sfix19_En18
  input [18:0] Wgt_0_246, // sfix19_En18
  input [18:0] Wgt_0_247, // sfix19_En18
  input [18:0] Wgt_0_248, // sfix19_En18
  input [18:0] Wgt_0_249, // sfix19_En18
  input [18:0] Wgt_0_250, // sfix19_En18
  input [18:0] Wgt_0_251, // sfix19_En18
  input [18:0] Wgt_0_252, // sfix19_En18
  input [18:0] Wgt_0_253, // sfix19_En18
  input [18:0] Wgt_0_254, // sfix19_En18
  input [18:0] Wgt_0_255, // sfix19_En18
  input [18:0] Wgt_0_256, // sfix19_En18
  input [18:0] Wgt_0_257, // sfix19_En18
  input [18:0] Wgt_0_258, // sfix19_En18
  input [18:0] Wgt_0_259, // sfix19_En18
  input [18:0] Wgt_0_260, // sfix19_En18
  input [18:0] Wgt_0_261, // sfix19_En18
  input [18:0] Wgt_0_262, // sfix19_En18
  input [18:0] Wgt_0_263, // sfix19_En18
  input [18:0] Wgt_0_264, // sfix19_En18
  input [18:0] Wgt_0_265, // sfix19_En18
  input [18:0] Wgt_0_266, // sfix19_En18
  input [18:0] Wgt_0_267, // sfix19_En18
  input [18:0] Wgt_0_268, // sfix19_En18
  input [18:0] Wgt_0_269, // sfix19_En18
  input [18:0] Wgt_0_270, // sfix19_En18
  input [18:0] Wgt_0_271, // sfix19_En18
  input [18:0] Wgt_0_272, // sfix19_En18
  input [18:0] Wgt_0_273, // sfix19_En18
  input [18:0] Wgt_0_274, // sfix19_En18
  input [18:0] Wgt_0_275, // sfix19_En18
  input [18:0] Wgt_0_276, // sfix19_En18
  input [18:0] Wgt_0_277, // sfix19_En18
  input [18:0] Wgt_0_278, // sfix19_En18
  input [18:0] Wgt_0_279, // sfix19_En18
  input [18:0] Wgt_0_280, // sfix19_En18
  input [18:0] Wgt_0_281, // sfix19_En18
  input [18:0] Wgt_0_282, // sfix19_En18
  input [18:0] Wgt_0_283, // sfix19_En18
  input [18:0] Wgt_0_284, // sfix19_En18
  input [18:0] Wgt_0_285, // sfix19_En18
  input [18:0] Wgt_0_286, // sfix19_En18
  input [18:0] Wgt_0_287, // sfix19_En18
  input [18:0] Wgt_0_288, // sfix19_En18
  input [18:0] Wgt_0_289, // sfix19_En18
  input [18:0] Wgt_0_290, // sfix19_En18
  input [18:0] Wgt_0_291, // sfix19_En18
  input [18:0] Wgt_0_292, // sfix19_En18
  input [18:0] Wgt_0_293, // sfix19_En18
  input [18:0] Wgt_0_294, // sfix19_En18
  input [18:0] Wgt_0_295, // sfix19_En18
  input [18:0] Wgt_0_296, // sfix19_En18
  input [18:0] Wgt_0_297, // sfix19_En18
  input [18:0] Wgt_0_298, // sfix19_En18
  input [18:0] Wgt_0_299, // sfix19_En18
  input [18:0] Wgt_0_300, // sfix19_En18
  input [18:0] Wgt_0_301, // sfix19_En18
  input [18:0] Wgt_0_302, // sfix19_En18
  input [18:0] Wgt_0_303, // sfix19_En18
  input [18:0] Wgt_0_304, // sfix19_En18
  input [18:0] Wgt_0_305, // sfix19_En18
  input [18:0] Wgt_0_306, // sfix19_En18
  input [18:0] Wgt_0_307, // sfix19_En18
  input [18:0] Wgt_0_308, // sfix19_En18
  input [18:0] Wgt_0_309, // sfix19_En18
  input [18:0] Wgt_0_310, // sfix19_En18
  input [18:0] Wgt_0_311, // sfix19_En18
  input [18:0] Wgt_0_312, // sfix19_En18
  input [18:0] Wgt_0_313, // sfix19_En18
  input [18:0] Wgt_0_314, // sfix19_En18
  input [18:0] Wgt_0_315, // sfix19_En18
  input [18:0] Wgt_0_316, // sfix19_En18
  input [18:0] Wgt_0_317, // sfix19_En18
  input [18:0] Wgt_0_318, // sfix19_En18
  input [18:0] Wgt_0_319, // sfix19_En18
  input [18:0] Wgt_0_320, // sfix19_En18
  input [18:0] Wgt_0_321, // sfix19_En18
  input [18:0] Wgt_0_322, // sfix19_En18
  input [18:0] Wgt_0_323, // sfix19_En18
  input [18:0] Wgt_0_324, // sfix19_En18
  input [18:0] Wgt_0_325, // sfix19_En18
  input [18:0] Wgt_0_326, // sfix19_En18
  input [18:0] Wgt_0_327, // sfix19_En18
  input [18:0] Wgt_0_328, // sfix19_En18
  input [18:0] Wgt_0_329, // sfix19_En18
  input [18:0] Wgt_0_330, // sfix19_En18
  input [18:0] Wgt_0_331, // sfix19_En18
  input [18:0] Wgt_0_332, // sfix19_En18
  input [18:0] Wgt_0_333, // sfix19_En18
  input [18:0] Wgt_0_334, // sfix19_En18
  input [18:0] Wgt_0_335, // sfix19_En18
  input [18:0] Wgt_0_336, // sfix19_En18
  input [18:0] Wgt_0_337, // sfix19_En18
  input [18:0] Wgt_0_338, // sfix19_En18
  input [18:0] Wgt_0_339, // sfix19_En18
  input [18:0] Wgt_0_340, // sfix19_En18
  input [18:0] Wgt_0_341, // sfix19_En18
  input [18:0] Wgt_0_342, // sfix19_En18
  input [18:0] Wgt_0_343, // sfix19_En18
  input [18:0] Wgt_0_344, // sfix19_En18
  input [18:0] Wgt_0_345, // sfix19_En18
  input [18:0] Wgt_0_346, // sfix19_En18
  input [18:0] Wgt_0_347, // sfix19_En18
  input [18:0] Wgt_0_348, // sfix19_En18
  input [18:0] Wgt_0_349, // sfix19_En18
  input [18:0] Wgt_0_350, // sfix19_En18
  input [18:0] Wgt_0_351, // sfix19_En18
  input [18:0] Wgt_0_352, // sfix19_En18
  input [18:0] Wgt_0_353, // sfix19_En18
  input [18:0] Wgt_0_354, // sfix19_En18
  input [18:0] Wgt_0_355, // sfix19_En18
  input [18:0] Wgt_0_356, // sfix19_En18
  input [18:0] Wgt_0_357, // sfix19_En18
  input [18:0] Wgt_0_358, // sfix19_En18
  input [18:0] Wgt_0_359, // sfix19_En18
  input [18:0] Wgt_0_360, // sfix19_En18
  input [18:0] Wgt_0_361, // sfix19_En18
  input [18:0] Wgt_0_362, // sfix19_En18
  input [18:0] Wgt_0_363, // sfix19_En18
  input [18:0] Wgt_0_364, // sfix19_En18
  input [18:0] Wgt_0_365, // sfix19_En18
  input [18:0] Wgt_0_366, // sfix19_En18
  input [18:0] Wgt_0_367, // sfix19_En18
  input [18:0] Wgt_0_368, // sfix19_En18
  input [18:0] Wgt_0_369, // sfix19_En18
  input [18:0] Wgt_0_370, // sfix19_En18
  input [18:0] Wgt_0_371, // sfix19_En18
  input [18:0] Wgt_0_372, // sfix19_En18
  input [18:0] Wgt_0_373, // sfix19_En18
  input [18:0] Wgt_0_374, // sfix19_En18
  input [18:0] Wgt_0_375, // sfix19_En18
  input [18:0] Wgt_0_376, // sfix19_En18
  input [18:0] Wgt_0_377, // sfix19_En18
  input [18:0] Wgt_0_378, // sfix19_En18
  input [18:0] Wgt_0_379, // sfix19_En18
  input [18:0] Wgt_0_380, // sfix19_En18
  input [18:0] Wgt_0_381, // sfix19_En18
  input [18:0] Wgt_0_382, // sfix19_En18
  input [18:0] Wgt_0_383, // sfix19_En18
  input [18:0] Wgt_0_384, // sfix19_En18
  input [18:0] Wgt_0_385, // sfix19_En18
  input [18:0] Wgt_0_386, // sfix19_En18
  input [18:0] Wgt_0_387, // sfix19_En18
  input [18:0] Wgt_0_388, // sfix19_En18
  input [18:0] Wgt_0_389, // sfix19_En18
  input [18:0] Wgt_0_390, // sfix19_En18
  input [18:0] Wgt_0_391, // sfix19_En18
  input [18:0] Wgt_0_392, // sfix19_En18
  input [18:0] Wgt_0_393, // sfix19_En18
  input [18:0] Wgt_0_394, // sfix19_En18
  input [18:0] Wgt_0_395, // sfix19_En18
  input [18:0] Wgt_0_396, // sfix19_En18
  input [18:0] Wgt_0_397, // sfix19_En18
  input [18:0] Wgt_0_398, // sfix19_En18
  input [18:0] Wgt_0_399, // sfix19_En18
  input [18:0] Wgt_0_400, // sfix19_En18
  input [18:0] Wgt_0_401, // sfix19_En18
  input [18:0] Wgt_0_402, // sfix19_En18
  input [18:0] Wgt_0_403, // sfix19_En18
  input [18:0] Wgt_0_404, // sfix19_En18
  input [18:0] Wgt_0_405, // sfix19_En18
  input [18:0] Wgt_0_406, // sfix19_En18
  input [18:0] Wgt_0_407, // sfix19_En18
  input [18:0] Wgt_0_408, // sfix19_En18
  input [18:0] Wgt_0_409, // sfix19_En18
  input [18:0] Wgt_0_410, // sfix19_En18
  input [18:0] Wgt_0_411, // sfix19_En18
  input [18:0] Wgt_0_412, // sfix19_En18
  input [18:0] Wgt_0_413, // sfix19_En18
  input [18:0] Wgt_0_414, // sfix19_En18
  input [18:0] Wgt_0_415, // sfix19_En18
  input [18:0] Wgt_0_416, // sfix19_En18
  input [18:0] Wgt_0_417, // sfix19_En18
  input [18:0] Wgt_0_418, // sfix19_En18
  input [18:0] Wgt_0_419, // sfix19_En18
  input [18:0] Wgt_0_420, // sfix19_En18
  input [18:0] Wgt_0_421, // sfix19_En18
  input [18:0] Wgt_0_422, // sfix19_En18
  input [18:0] Wgt_0_423, // sfix19_En18
  input [18:0] Wgt_0_424, // sfix19_En18
  input [18:0] Wgt_0_425, // sfix19_En18
  input [18:0] Wgt_0_426, // sfix19_En18
  input [18:0] Wgt_0_427, // sfix19_En18
  input [18:0] Wgt_0_428, // sfix19_En18
  input [18:0] Wgt_0_429, // sfix19_En18
  input [18:0] Wgt_0_430, // sfix19_En18
  input [18:0] Wgt_0_431, // sfix19_En18
  input [18:0] Wgt_0_432, // sfix19_En18
  input [18:0] Wgt_0_433, // sfix19_En18
  input [18:0] Wgt_0_434, // sfix19_En18
  input [18:0] Wgt_0_435, // sfix19_En18
  input [18:0] Wgt_0_436, // sfix19_En18
  input [18:0] Wgt_0_437, // sfix19_En18
  input [18:0] Wgt_0_438, // sfix19_En18
  input [18:0] Wgt_0_439, // sfix19_En18
  input [18:0] Wgt_0_440, // sfix19_En18
  input [18:0] Wgt_0_441, // sfix19_En18
  input [18:0] Wgt_0_442, // sfix19_En18
  input [18:0] Wgt_0_443, // sfix19_En18
  input [18:0] Wgt_0_444, // sfix19_En18
  input [18:0] Wgt_0_445, // sfix19_En18
  input [18:0] Wgt_0_446, // sfix19_En18
  input [18:0] Wgt_0_447, // sfix19_En18
  input [18:0] Wgt_0_448, // sfix19_En18
  input [18:0] Wgt_0_449, // sfix19_En18
  input [18:0] Wgt_0_450, // sfix19_En18
  input [18:0] Wgt_0_451, // sfix19_En18
  input [18:0] Wgt_0_452, // sfix19_En18
  input [18:0] Wgt_0_453, // sfix19_En18
  input [18:0] Wgt_0_454, // sfix19_En18
  input [18:0] Wgt_0_455, // sfix19_En18
  input [18:0] Wgt_0_456, // sfix19_En18
  input [18:0] Wgt_0_457, // sfix19_En18
  input [18:0] Wgt_0_458, // sfix19_En18
  input [18:0] Wgt_0_459, // sfix19_En18
  input [18:0] Wgt_0_460, // sfix19_En18
  input [18:0] Wgt_0_461, // sfix19_En18
  input [18:0] Wgt_0_462, // sfix19_En18
  input [18:0] Wgt_0_463, // sfix19_En18
  input [18:0] Wgt_0_464, // sfix19_En18
  input [18:0] Wgt_0_465, // sfix19_En18
  input [18:0] Wgt_0_466, // sfix19_En18
  input [18:0] Wgt_0_467, // sfix19_En18
  input [18:0] Wgt_0_468, // sfix19_En18
  input [18:0] Wgt_0_469, // sfix19_En18
  input [18:0] Wgt_0_470, // sfix19_En18
  input [18:0] Wgt_0_471, // sfix19_En18
  input [18:0] Wgt_0_472, // sfix19_En18
  input [18:0] Wgt_0_473, // sfix19_En18
  input [18:0] Wgt_0_474, // sfix19_En18
  input [18:0] Wgt_0_475, // sfix19_En18
  input [18:0] Wgt_0_476, // sfix19_En18
  input [18:0] Wgt_0_477, // sfix19_En18
  input [18:0] Wgt_0_478, // sfix19_En18
  input [18:0] Wgt_0_479, // sfix19_En18
  input [18:0] Wgt_0_480, // sfix19_En18
  input [18:0] Wgt_0_481, // sfix19_En18
  input [18:0] Wgt_0_482, // sfix19_En18
  input [18:0] Wgt_0_483, // sfix19_En18
  input [18:0] Wgt_0_484, // sfix19_En18
  input [18:0] Wgt_0_485, // sfix19_En18
  input [18:0] Wgt_0_486, // sfix19_En18
  input [18:0] Wgt_0_487, // sfix19_En18
  input [18:0] Wgt_0_488, // sfix19_En18
  input [18:0] Wgt_0_489, // sfix19_En18
  input [18:0] Wgt_0_490, // sfix19_En18
  input [18:0] Wgt_0_491, // sfix19_En18
  input [18:0] Wgt_0_492, // sfix19_En18
  input [18:0] Wgt_0_493, // sfix19_En18
  input [18:0] Wgt_0_494, // sfix19_En18
  input [18:0] Wgt_0_495, // sfix19_En18
  input [18:0] Wgt_0_496, // sfix19_En18
  input [18:0] Wgt_0_497, // sfix19_En18
  input [18:0] Wgt_0_498, // sfix19_En18
  input [18:0] Wgt_0_499, // sfix19_En18
  input [18:0] Wgt_0_500, // sfix19_En18
  input [18:0] Wgt_0_501, // sfix19_En18
  input [18:0] Wgt_0_502, // sfix19_En18
  input [18:0] Wgt_0_503, // sfix19_En18
  input [18:0] Wgt_0_504, // sfix19_En18
  input [18:0] Wgt_0_505, // sfix19_En18
  input [18:0] Wgt_0_506, // sfix19_En18
  input [18:0] Wgt_0_507, // sfix19_En18
  input [18:0] Wgt_0_508, // sfix19_En18
  input [18:0] Wgt_0_509, // sfix19_En18
  input [18:0] Wgt_0_510, // sfix19_En18
  input [18:0] Wgt_0_511, // sfix19_En18
  input [18:0] Wgt_0_512, // sfix19_En18
  input [18:0] Wgt_0_513, // sfix19_En18
  input [18:0] Wgt_0_514, // sfix19_En18
  input [18:0] Wgt_0_515, // sfix19_En18
  input [18:0] Wgt_0_516, // sfix19_En18
  input [18:0] Wgt_0_517, // sfix19_En18
  input [18:0] Wgt_0_518, // sfix19_En18
  input [18:0] Wgt_0_519, // sfix19_En18
  input [18:0] Wgt_0_520, // sfix19_En18
  input [18:0] Wgt_0_521, // sfix19_En18
  input [18:0] Wgt_0_522, // sfix19_En18
  input [18:0] Wgt_0_523, // sfix19_En18
  input [18:0] Wgt_0_524, // sfix19_En18
  input [18:0] Wgt_0_525, // sfix19_En18
  input [18:0] Wgt_0_526, // sfix19_En18
  input [18:0] Wgt_0_527, // sfix19_En18
  input [18:0] Wgt_0_528, // sfix19_En18
  input [18:0] Wgt_0_529, // sfix19_En18
  input [18:0] Wgt_0_530, // sfix19_En18
  input [18:0] Wgt_0_531, // sfix19_En18
  input [18:0] Wgt_0_532, // sfix19_En18
  input [18:0] Wgt_0_533, // sfix19_En18
  input [18:0] Wgt_0_534, // sfix19_En18
  input [18:0] Wgt_0_535, // sfix19_En18
  input [18:0] Wgt_0_536, // sfix19_En18
  input [18:0] Wgt_0_537, // sfix19_En18
  input [18:0] Wgt_0_538, // sfix19_En18
  input [18:0] Wgt_0_539, // sfix19_En18
  input [18:0] Wgt_0_540, // sfix19_En18
  input [18:0] Wgt_0_541, // sfix19_En18
  input [18:0] Wgt_0_542, // sfix19_En18
  input [18:0] Wgt_0_543, // sfix19_En18
  input [18:0] Wgt_0_544, // sfix19_En18
  input [18:0] Wgt_0_545, // sfix19_En18
  input [18:0] Wgt_0_546, // sfix19_En18
  input [18:0] Wgt_0_547, // sfix19_En18
  input [18:0] Wgt_0_548, // sfix19_En18
  input [18:0] Wgt_0_549, // sfix19_En18
  input [18:0] Wgt_0_550, // sfix19_En18
  input [18:0] Wgt_0_551, // sfix19_En18
  input [18:0] Wgt_0_552, // sfix19_En18
  input [18:0] Wgt_0_553, // sfix19_En18
  input [18:0] Wgt_0_554, // sfix19_En18
  input [18:0] Wgt_0_555, // sfix19_En18
  input [18:0] Wgt_0_556, // sfix19_En18
  input [18:0] Wgt_0_557, // sfix19_En18
  input [18:0] Wgt_0_558, // sfix19_En18
  input [18:0] Wgt_0_559, // sfix19_En18
  input [18:0] Wgt_0_560, // sfix19_En18
  input [18:0] Wgt_0_561, // sfix19_En18
  input [18:0] Wgt_0_562, // sfix19_En18
  input [18:0] Wgt_0_563, // sfix19_En18
  input [18:0] Wgt_0_564, // sfix19_En18
  input [18:0] Wgt_0_565, // sfix19_En18
  input [18:0] Wgt_0_566, // sfix19_En18
  input [18:0] Wgt_0_567, // sfix19_En18
  input [18:0] Wgt_0_568, // sfix19_En18
  input [18:0] Wgt_0_569, // sfix19_En18
  input [18:0] Wgt_0_570, // sfix19_En18
  input [18:0] Wgt_0_571, // sfix19_En18
  input [18:0] Wgt_0_572, // sfix19_En18
  input [18:0] Wgt_0_573, // sfix19_En18
  input [18:0] Wgt_0_574, // sfix19_En18
  input [18:0] Wgt_0_575, // sfix19_En18
  input [18:0] Wgt_0_576, // sfix19_En18
  input [18:0] Wgt_0_577, // sfix19_En18
  input [18:0] Wgt_0_578, // sfix19_En18
  input [18:0] Wgt_0_579, // sfix19_En18
  input [18:0] Wgt_0_580, // sfix19_En18
  input [18:0] Wgt_0_581, // sfix19_En18
  input [18:0] Wgt_0_582, // sfix19_En18
  input [18:0] Wgt_0_583, // sfix19_En18
  input [18:0] Wgt_0_584, // sfix19_En18
  input [18:0] Wgt_0_585, // sfix19_En18
  input [18:0] Wgt_0_586, // sfix19_En18
  input [18:0] Wgt_0_587, // sfix19_En18
  input [18:0] Wgt_0_588, // sfix19_En18
  input [18:0] Wgt_0_589, // sfix19_En18
  input [18:0] Wgt_0_590, // sfix19_En18
  input [18:0] Wgt_0_591, // sfix19_En18
  input [18:0] Wgt_0_592, // sfix19_En18
  input [18:0] Wgt_0_593, // sfix19_En18
  input [18:0] Wgt_0_594, // sfix19_En18
  input [18:0] Wgt_0_595, // sfix19_En18
  input [18:0] Wgt_0_596, // sfix19_En18
  input [18:0] Wgt_0_597, // sfix19_En18
  input [18:0] Wgt_0_598, // sfix19_En18
  input [18:0] Wgt_0_599, // sfix19_En18
  input [18:0] Wgt_0_600, // sfix19_En18
  input [18:0] Wgt_0_601, // sfix19_En18
  input [18:0] Wgt_0_602, // sfix19_En18
  input [18:0] Wgt_0_603, // sfix19_En18
  input [18:0] Wgt_0_604, // sfix19_En18
  input [18:0] Wgt_0_605, // sfix19_En18
  input [18:0] Wgt_0_606, // sfix19_En18
  input [18:0] Wgt_0_607, // sfix19_En18
  input [18:0] Wgt_0_608, // sfix19_En18
  input [18:0] Wgt_0_609, // sfix19_En18
  input [18:0] Wgt_0_610, // sfix19_En18
  input [18:0] Wgt_0_611, // sfix19_En18
  input [18:0] Wgt_0_612, // sfix19_En18
  input [18:0] Wgt_0_613, // sfix19_En18
  input [18:0] Wgt_0_614, // sfix19_En18
  input [18:0] Wgt_0_615, // sfix19_En18
  input [18:0] Wgt_0_616, // sfix19_En18
  input [18:0] Wgt_0_617, // sfix19_En18
  input [18:0] Wgt_0_618, // sfix19_En18
  input [18:0] Wgt_0_619, // sfix19_En18
  input [18:0] Wgt_0_620, // sfix19_En18
  input [18:0] Wgt_0_621, // sfix19_En18
  input [18:0] Wgt_0_622, // sfix19_En18
  input [18:0] Wgt_0_623, // sfix19_En18
  input [18:0] Wgt_0_624, // sfix19_En18
  input [18:0] Wgt_0_625, // sfix19_En18
  input [18:0] Wgt_0_626, // sfix19_En18
  input [18:0] Wgt_0_627, // sfix19_En18
  input [18:0] Wgt_0_628, // sfix19_En18
  input [18:0] Wgt_0_629, // sfix19_En18
  input [18:0] Wgt_0_630, // sfix19_En18
  input [18:0] Wgt_0_631, // sfix19_En18
  input [18:0] Wgt_0_632, // sfix19_En18
  input [18:0] Wgt_0_633, // sfix19_En18
  input [18:0] Wgt_0_634, // sfix19_En18
  input [18:0] Wgt_0_635, // sfix19_En18
  input [18:0] Wgt_0_636, // sfix19_En18
  input [18:0] Wgt_0_637, // sfix19_En18
  input [18:0] Wgt_0_638, // sfix19_En18
  input [18:0] Wgt_0_639, // sfix19_En18
  input [18:0] Wgt_0_640, // sfix19_En18
  input [18:0] Wgt_0_641, // sfix19_En18
  input [18:0] Wgt_0_642, // sfix19_En18
  input [18:0] Wgt_0_643, // sfix19_En18
  input [18:0] Wgt_0_644, // sfix19_En18
  input [18:0] Wgt_0_645, // sfix19_En18
  input [18:0] Wgt_0_646, // sfix19_En18
  input [18:0] Wgt_0_647, // sfix19_En18
  input [18:0] Wgt_0_648, // sfix19_En18
  input [18:0] Wgt_0_649, // sfix19_En18
  input [18:0] Wgt_0_650, // sfix19_En18
  input [18:0] Wgt_0_651, // sfix19_En18
  input [18:0] Wgt_0_652, // sfix19_En18
  input [18:0] Wgt_0_653, // sfix19_En18
  input [18:0] Wgt_0_654, // sfix19_En18
  input [18:0] Wgt_0_655, // sfix19_En18
  input [18:0] Wgt_0_656, // sfix19_En18
  input [18:0] Wgt_0_657, // sfix19_En18
  input [18:0] Wgt_0_658, // sfix19_En18
  input [18:0] Wgt_0_659, // sfix19_En18
  input [18:0] Wgt_0_660, // sfix19_En18
  input [18:0] Wgt_0_661, // sfix19_En18
  input [18:0] Wgt_0_662, // sfix19_En18
  input [18:0] Wgt_0_663, // sfix19_En18
  input [18:0] Wgt_0_664, // sfix19_En18
  input [18:0] Wgt_0_665, // sfix19_En18
  input [18:0] Wgt_0_666, // sfix19_En18
  input [18:0] Wgt_0_667, // sfix19_En18
  input [18:0] Wgt_0_668, // sfix19_En18
  input [18:0] Wgt_0_669, // sfix19_En18
  input [18:0] Wgt_0_670, // sfix19_En18
  input [18:0] Wgt_0_671, // sfix19_En18
  input [18:0] Wgt_0_672, // sfix19_En18
  input [18:0] Wgt_0_673, // sfix19_En18
  input [18:0] Wgt_0_674, // sfix19_En18
  input [18:0] Wgt_0_675, // sfix19_En18
  input [18:0] Wgt_0_676, // sfix19_En18
  input [18:0] Wgt_0_677, // sfix19_En18
  input [18:0] Wgt_0_678, // sfix19_En18
  input [18:0] Wgt_0_679, // sfix19_En18
  input [18:0] Wgt_0_680, // sfix19_En18
  input [18:0] Wgt_0_681, // sfix19_En18
  input [18:0] Wgt_0_682, // sfix19_En18
  input [18:0] Wgt_0_683, // sfix19_En18
  input [18:0] Wgt_0_684, // sfix19_En18
  input [18:0] Wgt_0_685, // sfix19_En18
  input [18:0] Wgt_0_686, // sfix19_En18
  input [18:0] Wgt_0_687, // sfix19_En18
  input [18:0] Wgt_0_688, // sfix19_En18
  input [18:0] Wgt_0_689, // sfix19_En18
  input [18:0] Wgt_0_690, // sfix19_En18
  input [18:0] Wgt_0_691, // sfix19_En18
  input [18:0] Wgt_0_692, // sfix19_En18
  input [18:0] Wgt_0_693, // sfix19_En18
  input [18:0] Wgt_0_694, // sfix19_En18
  input [18:0] Wgt_0_695, // sfix19_En18
  input [18:0] Wgt_0_696, // sfix19_En18
  input [18:0] Wgt_0_697, // sfix19_En18
  input [18:0] Wgt_0_698, // sfix19_En18
  input [18:0] Wgt_0_699, // sfix19_En18
  input [18:0] Wgt_0_700, // sfix19_En18
  input [18:0] Wgt_0_701, // sfix19_En18
  input [18:0] Wgt_0_702, // sfix19_En18
  input [18:0] Wgt_0_703, // sfix19_En18
  input [18:0] Wgt_0_704, // sfix19_En18
  input [18:0] Wgt_0_705, // sfix19_En18
  input [18:0] Wgt_0_706, // sfix19_En18
  input [18:0] Wgt_0_707, // sfix19_En18
  input [18:0] Wgt_0_708, // sfix19_En18
  input [18:0] Wgt_0_709, // sfix19_En18
  input [18:0] Wgt_0_710, // sfix19_En18
  input [18:0] Wgt_0_711, // sfix19_En18
  input [18:0] Wgt_0_712, // sfix19_En18
  input [18:0] Wgt_0_713, // sfix19_En18
  input [18:0] Wgt_0_714, // sfix19_En18
  input [18:0] Wgt_0_715, // sfix19_En18
  input [18:0] Wgt_0_716, // sfix19_En18
  input [18:0] Wgt_0_717, // sfix19_En18
  input [18:0] Wgt_0_718, // sfix19_En18
  input [18:0] Wgt_0_719, // sfix19_En18
  input [18:0] Wgt_0_720, // sfix19_En18
  input [18:0] Wgt_0_721, // sfix19_En18
  input [18:0] Wgt_0_722, // sfix19_En18
  input [18:0] Wgt_0_723, // sfix19_En18
  input [18:0] Wgt_0_724, // sfix19_En18
  input [18:0] Wgt_0_725, // sfix19_En18
  input [18:0] Wgt_0_726, // sfix19_En18
  input [18:0] Wgt_0_727, // sfix19_En18
  input [18:0] Wgt_0_728, // sfix19_En18
  input [18:0] Wgt_0_729, // sfix19_En18
  input [18:0] Wgt_0_730, // sfix19_En18
  input [18:0] Wgt_0_731, // sfix19_En18
  input [18:0] Wgt_0_732, // sfix19_En18
  input [18:0] Wgt_0_733, // sfix19_En18
  input [18:0] Wgt_0_734, // sfix19_En18
  input [18:0] Wgt_0_735, // sfix19_En18
  input [18:0] Wgt_0_736, // sfix19_En18
  input [18:0] Wgt_0_737, // sfix19_En18
  input [18:0] Wgt_0_738, // sfix19_En18
  input [18:0] Wgt_0_739, // sfix19_En18
  input [18:0] Wgt_0_740, // sfix19_En18
  input [18:0] Wgt_0_741, // sfix19_En18
  input [18:0] Wgt_0_742, // sfix19_En18
  input [18:0] Wgt_0_743, // sfix19_En18
  input [18:0] Wgt_0_744, // sfix19_En18
  input [18:0] Wgt_0_745, // sfix19_En18
  input [18:0] Wgt_0_746, // sfix19_En18
  input [18:0] Wgt_0_747, // sfix19_En18
  input [18:0] Wgt_0_748, // sfix19_En18
  input [18:0] Wgt_0_749, // sfix19_En18
  input [18:0] Wgt_0_750, // sfix19_En18
  input [18:0] Wgt_0_751, // sfix19_En18
  input [18:0] Wgt_0_752, // sfix19_En18
  input [18:0] Wgt_0_753, // sfix19_En18
  input [18:0] Wgt_0_754, // sfix19_En18
  input [18:0] Wgt_0_755, // sfix19_En18
  input [18:0] Wgt_0_756, // sfix19_En18
  input [18:0] Wgt_0_757, // sfix19_En18
  input [18:0] Wgt_0_758, // sfix19_En18
  input [18:0] Wgt_0_759, // sfix19_En18
  input [18:0] Wgt_0_760, // sfix19_En18
  input [18:0] Wgt_0_761, // sfix19_En18
  input [18:0] Wgt_0_762, // sfix19_En18
  input [18:0] Wgt_0_763, // sfix19_En18
  input [18:0] Wgt_0_764, // sfix19_En18
  input [18:0] Wgt_0_765, // sfix19_En18
  input [18:0] Wgt_0_766, // sfix19_En18
  input [18:0] Wgt_0_767, // sfix19_En18
  input [18:0] Wgt_0_768, // sfix19_En18
  input [18:0] Wgt_0_769, // sfix19_En18
  input [18:0] Wgt_0_770, // sfix19_En18
  input [18:0] Wgt_0_771, // sfix19_En18
  input [18:0] Wgt_0_772, // sfix19_En18
  input [18:0] Wgt_0_773, // sfix19_En18
  input [18:0] Wgt_0_774, // sfix19_En18
  input [18:0] Wgt_0_775, // sfix19_En18
  input [18:0] Wgt_0_776, // sfix19_En18
  input [18:0] Wgt_0_777, // sfix19_En18
  input [18:0] Wgt_0_778, // sfix19_En18
  input [18:0] Wgt_0_779, // sfix19_En18
  input [18:0] Wgt_0_780, // sfix19_En18
  input [18:0] Wgt_0_781, // sfix19_En18
  input [18:0] Wgt_0_782, // sfix19_En18
  input [18:0] Wgt_0_783, // sfix19_En18
  input [18:0] Wgt_0_784, // sfix19_En18
  input [18:0] Wgt_1_0, // sfix19_En18
  input [18:0] Wgt_1_1, // sfix19_En18
  input [18:0] Wgt_1_2, // sfix19_En18
  input [18:0] Wgt_1_3, // sfix19_En18
  input [18:0] Wgt_1_4, // sfix19_En18
  input [18:0] Wgt_1_5, // sfix19_En18
  input [18:0] Wgt_1_6, // sfix19_En18
  input [18:0] Wgt_1_7, // sfix19_En18
  input [18:0] Wgt_1_8, // sfix19_En18
  input [18:0] Wgt_1_9, // sfix19_En18
  input [18:0] Wgt_1_10, // sfix19_En18
  input [18:0] Wgt_1_11, // sfix19_En18
  input [18:0] Wgt_1_12, // sfix19_En18
  input [18:0] Wgt_1_13, // sfix19_En18
  input [18:0] Wgt_1_14, // sfix19_En18
  input [18:0] Wgt_1_15, // sfix19_En18
  input [18:0] Wgt_1_16, // sfix19_En18
  input [18:0] Wgt_1_17, // sfix19_En18
  input [18:0] Wgt_1_18, // sfix19_En18
  input [18:0] Wgt_1_19, // sfix19_En18
  input [18:0] Wgt_1_20, // sfix19_En18
  input [18:0] Wgt_1_21, // sfix19_En18
  input [18:0] Wgt_1_22, // sfix19_En18
  input [18:0] Wgt_1_23, // sfix19_En18
  input [18:0] Wgt_1_24, // sfix19_En18
  input [18:0] Wgt_1_25, // sfix19_En18
  input [18:0] Wgt_1_26, // sfix19_En18
  input [18:0] Wgt_1_27, // sfix19_En18
  input [18:0] Wgt_1_28, // sfix19_En18
  input [18:0] Wgt_1_29, // sfix19_En18
  input [18:0] Wgt_1_30, // sfix19_En18
  input [18:0] Wgt_1_31, // sfix19_En18
  input [18:0] Wgt_1_32, // sfix19_En18
  input [18:0] Wgt_1_33, // sfix19_En18
  input [18:0] Wgt_1_34, // sfix19_En18
  input [18:0] Wgt_1_35, // sfix19_En18
  input [18:0] Wgt_1_36, // sfix19_En18
  input [18:0] Wgt_1_37, // sfix19_En18
  input [18:0] Wgt_1_38, // sfix19_En18
  input [18:0] Wgt_1_39, // sfix19_En18
  input [18:0] Wgt_1_40, // sfix19_En18
  input [18:0] Wgt_1_41, // sfix19_En18
  input [18:0] Wgt_1_42, // sfix19_En18
  input [18:0] Wgt_1_43, // sfix19_En18
  input [18:0] Wgt_1_44, // sfix19_En18
  input [18:0] Wgt_1_45, // sfix19_En18
  input [18:0] Wgt_1_46, // sfix19_En18
  input [18:0] Wgt_1_47, // sfix19_En18
  input [18:0] Wgt_1_48, // sfix19_En18
  input [18:0] Wgt_1_49, // sfix19_En18
  input [18:0] Wgt_1_50, // sfix19_En18
  input [18:0] Wgt_1_51, // sfix19_En18
  input [18:0] Wgt_1_52, // sfix19_En18
  input [18:0] Wgt_1_53, // sfix19_En18
  input [18:0] Wgt_1_54, // sfix19_En18
  input [18:0] Wgt_1_55, // sfix19_En18
  input [18:0] Wgt_1_56, // sfix19_En18
  input [18:0] Wgt_1_57, // sfix19_En18
  input [18:0] Wgt_1_58, // sfix19_En18
  input [18:0] Wgt_1_59, // sfix19_En18
  input [18:0] Wgt_1_60, // sfix19_En18
  input [18:0] Wgt_1_61, // sfix19_En18
  input [18:0] Wgt_1_62, // sfix19_En18
  input [18:0] Wgt_1_63, // sfix19_En18
  input [18:0] Wgt_1_64, // sfix19_En18
  input [18:0] Wgt_1_65, // sfix19_En18
  input [18:0] Wgt_1_66, // sfix19_En18
  input [18:0] Wgt_1_67, // sfix19_En18
  input [18:0] Wgt_1_68, // sfix19_En18
  input [18:0] Wgt_1_69, // sfix19_En18
  input [18:0] Wgt_1_70, // sfix19_En18
  input [18:0] Wgt_1_71, // sfix19_En18
  input [18:0] Wgt_1_72, // sfix19_En18
  input [18:0] Wgt_1_73, // sfix19_En18
  input [18:0] Wgt_1_74, // sfix19_En18
  input [18:0] Wgt_1_75, // sfix19_En18
  input [18:0] Wgt_1_76, // sfix19_En18
  input [18:0] Wgt_1_77, // sfix19_En18
  input [18:0] Wgt_1_78, // sfix19_En18
  input [18:0] Wgt_1_79, // sfix19_En18
  input [18:0] Wgt_1_80, // sfix19_En18
  input [18:0] Wgt_1_81, // sfix19_En18
  input [18:0] Wgt_1_82, // sfix19_En18
  input [18:0] Wgt_1_83, // sfix19_En18
  input [18:0] Wgt_1_84, // sfix19_En18
  input [18:0] Wgt_1_85, // sfix19_En18
  input [18:0] Wgt_1_86, // sfix19_En18
  input [18:0] Wgt_1_87, // sfix19_En18
  input [18:0] Wgt_1_88, // sfix19_En18
  input [18:0] Wgt_1_89, // sfix19_En18
  input [18:0] Wgt_1_90, // sfix19_En18
  input [18:0] Wgt_1_91, // sfix19_En18
  input [18:0] Wgt_1_92, // sfix19_En18
  input [18:0] Wgt_1_93, // sfix19_En18
  input [18:0] Wgt_1_94, // sfix19_En18
  input [18:0] Wgt_1_95, // sfix19_En18
  input [18:0] Wgt_1_96, // sfix19_En18
  input [18:0] Wgt_1_97, // sfix19_En18
  input [18:0] Wgt_1_98, // sfix19_En18
  input [18:0] Wgt_1_99, // sfix19_En18
  input [18:0] Wgt_1_100, // sfix19_En18
  input [18:0] Wgt_1_101, // sfix19_En18
  input [18:0] Wgt_1_102, // sfix19_En18
  input [18:0] Wgt_1_103, // sfix19_En18
  input [18:0] Wgt_1_104, // sfix19_En18
  input [18:0] Wgt_1_105, // sfix19_En18
  input [18:0] Wgt_1_106, // sfix19_En18
  input [18:0] Wgt_1_107, // sfix19_En18
  input [18:0] Wgt_1_108, // sfix19_En18
  input [18:0] Wgt_1_109, // sfix19_En18
  input [18:0] Wgt_1_110, // sfix19_En18
  input [18:0] Wgt_1_111, // sfix19_En18
  input [18:0] Wgt_1_112, // sfix19_En18
  input [18:0] Wgt_1_113, // sfix19_En18
  input [18:0] Wgt_1_114, // sfix19_En18
  input [18:0] Wgt_1_115, // sfix19_En18
  input [18:0] Wgt_1_116, // sfix19_En18
  input [18:0] Wgt_1_117, // sfix19_En18
  input [18:0] Wgt_1_118, // sfix19_En18
  input [18:0] Wgt_1_119, // sfix19_En18
  input [18:0] Wgt_1_120, // sfix19_En18
  input [18:0] Wgt_1_121, // sfix19_En18
  input [18:0] Wgt_1_122, // sfix19_En18
  input [18:0] Wgt_1_123, // sfix19_En18
  input [18:0] Wgt_1_124, // sfix19_En18
  input [18:0] Wgt_1_125, // sfix19_En18
  input [18:0] Wgt_1_126, // sfix19_En18
  input [18:0] Wgt_1_127, // sfix19_En18
  input [18:0] Wgt_1_128, // sfix19_En18
  input [18:0] Wgt_1_129, // sfix19_En18
  input [18:0] Wgt_1_130, // sfix19_En18
  input [18:0] Wgt_1_131, // sfix19_En18
  input [18:0] Wgt_1_132, // sfix19_En18
  input [18:0] Wgt_1_133, // sfix19_En18
  input [18:0] Wgt_1_134, // sfix19_En18
  input [18:0] Wgt_1_135, // sfix19_En18
  input [18:0] Wgt_1_136, // sfix19_En18
  input [18:0] Wgt_1_137, // sfix19_En18
  input [18:0] Wgt_1_138, // sfix19_En18
  input [18:0] Wgt_1_139, // sfix19_En18
  input [18:0] Wgt_1_140, // sfix19_En18
  input [18:0] Wgt_1_141, // sfix19_En18
  input [18:0] Wgt_1_142, // sfix19_En18
  input [18:0] Wgt_1_143, // sfix19_En18
  input [18:0] Wgt_1_144, // sfix19_En18
  input [18:0] Wgt_1_145, // sfix19_En18
  input [18:0] Wgt_1_146, // sfix19_En18
  input [18:0] Wgt_1_147, // sfix19_En18
  input [18:0] Wgt_1_148, // sfix19_En18
  input [18:0] Wgt_1_149, // sfix19_En18
  input [18:0] Wgt_1_150, // sfix19_En18
  input [18:0] Wgt_1_151, // sfix19_En18
  input [18:0] Wgt_1_152, // sfix19_En18
  input [18:0] Wgt_1_153, // sfix19_En18
  input [18:0] Wgt_1_154, // sfix19_En18
  input [18:0] Wgt_1_155, // sfix19_En18
  input [18:0] Wgt_1_156, // sfix19_En18
  input [18:0] Wgt_1_157, // sfix19_En18
  input [18:0] Wgt_1_158, // sfix19_En18
  input [18:0] Wgt_1_159, // sfix19_En18
  input [18:0] Wgt_1_160, // sfix19_En18
  input [18:0] Wgt_1_161, // sfix19_En18
  input [18:0] Wgt_1_162, // sfix19_En18
  input [18:0] Wgt_1_163, // sfix19_En18
  input [18:0] Wgt_1_164, // sfix19_En18
  input [18:0] Wgt_1_165, // sfix19_En18
  input [18:0] Wgt_1_166, // sfix19_En18
  input [18:0] Wgt_1_167, // sfix19_En18
  input [18:0] Wgt_1_168, // sfix19_En18
  input [18:0] Wgt_1_169, // sfix19_En18
  input [18:0] Wgt_1_170, // sfix19_En18
  input [18:0] Wgt_1_171, // sfix19_En18
  input [18:0] Wgt_1_172, // sfix19_En18
  input [18:0] Wgt_1_173, // sfix19_En18
  input [18:0] Wgt_1_174, // sfix19_En18
  input [18:0] Wgt_1_175, // sfix19_En18
  input [18:0] Wgt_1_176, // sfix19_En18
  input [18:0] Wgt_1_177, // sfix19_En18
  input [18:0] Wgt_1_178, // sfix19_En18
  input [18:0] Wgt_1_179, // sfix19_En18
  input [18:0] Wgt_1_180, // sfix19_En18
  input [18:0] Wgt_1_181, // sfix19_En18
  input [18:0] Wgt_1_182, // sfix19_En18
  input [18:0] Wgt_1_183, // sfix19_En18
  input [18:0] Wgt_1_184, // sfix19_En18
  input [18:0] Wgt_1_185, // sfix19_En18
  input [18:0] Wgt_1_186, // sfix19_En18
  input [18:0] Wgt_1_187, // sfix19_En18
  input [18:0] Wgt_1_188, // sfix19_En18
  input [18:0] Wgt_1_189, // sfix19_En18
  input [18:0] Wgt_1_190, // sfix19_En18
  input [18:0] Wgt_1_191, // sfix19_En18
  input [18:0] Wgt_1_192, // sfix19_En18
  input [18:0] Wgt_1_193, // sfix19_En18
  input [18:0] Wgt_1_194, // sfix19_En18
  input [18:0] Wgt_1_195, // sfix19_En18
  input [18:0] Wgt_1_196, // sfix19_En18
  input [18:0] Wgt_1_197, // sfix19_En18
  input [18:0] Wgt_1_198, // sfix19_En18
  input [18:0] Wgt_1_199, // sfix19_En18
  input [18:0] Wgt_1_200, // sfix19_En18
  input [18:0] Wgt_1_201, // sfix19_En18
  input [18:0] Wgt_1_202, // sfix19_En18
  input [18:0] Wgt_1_203, // sfix19_En18
  input [18:0] Wgt_1_204, // sfix19_En18
  input [18:0] Wgt_1_205, // sfix19_En18
  input [18:0] Wgt_1_206, // sfix19_En18
  input [18:0] Wgt_1_207, // sfix19_En18
  input [18:0] Wgt_1_208, // sfix19_En18
  input [18:0] Wgt_1_209, // sfix19_En18
  input [18:0] Wgt_1_210, // sfix19_En18
  input [18:0] Wgt_1_211, // sfix19_En18
  input [18:0] Wgt_1_212, // sfix19_En18
  input [18:0] Wgt_1_213, // sfix19_En18
  input [18:0] Wgt_1_214, // sfix19_En18
  input [18:0] Wgt_1_215, // sfix19_En18
  input [18:0] Wgt_1_216, // sfix19_En18
  input [18:0] Wgt_1_217, // sfix19_En18
  input [18:0] Wgt_1_218, // sfix19_En18
  input [18:0] Wgt_1_219, // sfix19_En18
  input [18:0] Wgt_1_220, // sfix19_En18
  input [18:0] Wgt_1_221, // sfix19_En18
  input [18:0] Wgt_1_222, // sfix19_En18
  input [18:0] Wgt_1_223, // sfix19_En18
  input [18:0] Wgt_1_224, // sfix19_En18
  input [18:0] Wgt_1_225, // sfix19_En18
  input [18:0] Wgt_1_226, // sfix19_En18
  input [18:0] Wgt_1_227, // sfix19_En18
  input [18:0] Wgt_1_228, // sfix19_En18
  input [18:0] Wgt_1_229, // sfix19_En18
  input [18:0] Wgt_1_230, // sfix19_En18
  input [18:0] Wgt_1_231, // sfix19_En18
  input [18:0] Wgt_1_232, // sfix19_En18
  input [18:0] Wgt_1_233, // sfix19_En18
  input [18:0] Wgt_1_234, // sfix19_En18
  input [18:0] Wgt_1_235, // sfix19_En18
  input [18:0] Wgt_1_236, // sfix19_En18
  input [18:0] Wgt_1_237, // sfix19_En18
  input [18:0] Wgt_1_238, // sfix19_En18
  input [18:0] Wgt_1_239, // sfix19_En18
  input [18:0] Wgt_1_240, // sfix19_En18
  input [18:0] Wgt_1_241, // sfix19_En18
  input [18:0] Wgt_1_242, // sfix19_En18
  input [18:0] Wgt_1_243, // sfix19_En18
  input [18:0] Wgt_1_244, // sfix19_En18
  input [18:0] Wgt_1_245, // sfix19_En18
  input [18:0] Wgt_1_246, // sfix19_En18
  input [18:0] Wgt_1_247, // sfix19_En18
  input [18:0] Wgt_1_248, // sfix19_En18
  input [18:0] Wgt_1_249, // sfix19_En18
  input [18:0] Wgt_1_250, // sfix19_En18
  input [18:0] Wgt_1_251, // sfix19_En18
  input [18:0] Wgt_1_252, // sfix19_En18
  input [18:0] Wgt_1_253, // sfix19_En18
  input [18:0] Wgt_1_254, // sfix19_En18
  input [18:0] Wgt_1_255, // sfix19_En18
  input [18:0] Wgt_1_256, // sfix19_En18
  input [18:0] Wgt_1_257, // sfix19_En18
  input [18:0] Wgt_1_258, // sfix19_En18
  input [18:0] Wgt_1_259, // sfix19_En18
  input [18:0] Wgt_1_260, // sfix19_En18
  input [18:0] Wgt_1_261, // sfix19_En18
  input [18:0] Wgt_1_262, // sfix19_En18
  input [18:0] Wgt_1_263, // sfix19_En18
  input [18:0] Wgt_1_264, // sfix19_En18
  input [18:0] Wgt_1_265, // sfix19_En18
  input [18:0] Wgt_1_266, // sfix19_En18
  input [18:0] Wgt_1_267, // sfix19_En18
  input [18:0] Wgt_1_268, // sfix19_En18
  input [18:0] Wgt_1_269, // sfix19_En18
  input [18:0] Wgt_1_270, // sfix19_En18
  input [18:0] Wgt_1_271, // sfix19_En18
  input [18:0] Wgt_1_272, // sfix19_En18
  input [18:0] Wgt_1_273, // sfix19_En18
  input [18:0] Wgt_1_274, // sfix19_En18
  input [18:0] Wgt_1_275, // sfix19_En18
  input [18:0] Wgt_1_276, // sfix19_En18
  input [18:0] Wgt_1_277, // sfix19_En18
  input [18:0] Wgt_1_278, // sfix19_En18
  input [18:0] Wgt_1_279, // sfix19_En18
  input [18:0] Wgt_1_280, // sfix19_En18
  input [18:0] Wgt_1_281, // sfix19_En18
  input [18:0] Wgt_1_282, // sfix19_En18
  input [18:0] Wgt_1_283, // sfix19_En18
  input [18:0] Wgt_1_284, // sfix19_En18
  input [18:0] Wgt_1_285, // sfix19_En18
  input [18:0] Wgt_1_286, // sfix19_En18
  input [18:0] Wgt_1_287, // sfix19_En18
  input [18:0] Wgt_1_288, // sfix19_En18
  input [18:0] Wgt_1_289, // sfix19_En18
  input [18:0] Wgt_1_290, // sfix19_En18
  input [18:0] Wgt_1_291, // sfix19_En18
  input [18:0] Wgt_1_292, // sfix19_En18
  input [18:0] Wgt_1_293, // sfix19_En18
  input [18:0] Wgt_1_294, // sfix19_En18
  input [18:0] Wgt_1_295, // sfix19_En18
  input [18:0] Wgt_1_296, // sfix19_En18
  input [18:0] Wgt_1_297, // sfix19_En18
  input [18:0] Wgt_1_298, // sfix19_En18
  input [18:0] Wgt_1_299, // sfix19_En18
  input [18:0] Wgt_1_300, // sfix19_En18
  input [18:0] Wgt_1_301, // sfix19_En18
  input [18:0] Wgt_1_302, // sfix19_En18
  input [18:0] Wgt_1_303, // sfix19_En18
  input [18:0] Wgt_1_304, // sfix19_En18
  input [18:0] Wgt_1_305, // sfix19_En18
  input [18:0] Wgt_1_306, // sfix19_En18
  input [18:0] Wgt_1_307, // sfix19_En18
  input [18:0] Wgt_1_308, // sfix19_En18
  input [18:0] Wgt_1_309, // sfix19_En18
  input [18:0] Wgt_1_310, // sfix19_En18
  input [18:0] Wgt_1_311, // sfix19_En18
  input [18:0] Wgt_1_312, // sfix19_En18
  input [18:0] Wgt_1_313, // sfix19_En18
  input [18:0] Wgt_1_314, // sfix19_En18
  input [18:0] Wgt_1_315, // sfix19_En18
  input [18:0] Wgt_1_316, // sfix19_En18
  input [18:0] Wgt_1_317, // sfix19_En18
  input [18:0] Wgt_1_318, // sfix19_En18
  input [18:0] Wgt_1_319, // sfix19_En18
  input [18:0] Wgt_1_320, // sfix19_En18
  input [18:0] Wgt_1_321, // sfix19_En18
  input [18:0] Wgt_1_322, // sfix19_En18
  input [18:0] Wgt_1_323, // sfix19_En18
  input [18:0] Wgt_1_324, // sfix19_En18
  input [18:0] Wgt_1_325, // sfix19_En18
  input [18:0] Wgt_1_326, // sfix19_En18
  input [18:0] Wgt_1_327, // sfix19_En18
  input [18:0] Wgt_1_328, // sfix19_En18
  input [18:0] Wgt_1_329, // sfix19_En18
  input [18:0] Wgt_1_330, // sfix19_En18
  input [18:0] Wgt_1_331, // sfix19_En18
  input [18:0] Wgt_1_332, // sfix19_En18
  input [18:0] Wgt_1_333, // sfix19_En18
  input [18:0] Wgt_1_334, // sfix19_En18
  input [18:0] Wgt_1_335, // sfix19_En18
  input [18:0] Wgt_1_336, // sfix19_En18
  input [18:0] Wgt_1_337, // sfix19_En18
  input [18:0] Wgt_1_338, // sfix19_En18
  input [18:0] Wgt_1_339, // sfix19_En18
  input [18:0] Wgt_1_340, // sfix19_En18
  input [18:0] Wgt_1_341, // sfix19_En18
  input [18:0] Wgt_1_342, // sfix19_En18
  input [18:0] Wgt_1_343, // sfix19_En18
  input [18:0] Wgt_1_344, // sfix19_En18
  input [18:0] Wgt_1_345, // sfix19_En18
  input [18:0] Wgt_1_346, // sfix19_En18
  input [18:0] Wgt_1_347, // sfix19_En18
  input [18:0] Wgt_1_348, // sfix19_En18
  input [18:0] Wgt_1_349, // sfix19_En18
  input [18:0] Wgt_1_350, // sfix19_En18
  input [18:0] Wgt_1_351, // sfix19_En18
  input [18:0] Wgt_1_352, // sfix19_En18
  input [18:0] Wgt_1_353, // sfix19_En18
  input [18:0] Wgt_1_354, // sfix19_En18
  input [18:0] Wgt_1_355, // sfix19_En18
  input [18:0] Wgt_1_356, // sfix19_En18
  input [18:0] Wgt_1_357, // sfix19_En18
  input [18:0] Wgt_1_358, // sfix19_En18
  input [18:0] Wgt_1_359, // sfix19_En18
  input [18:0] Wgt_1_360, // sfix19_En18
  input [18:0] Wgt_1_361, // sfix19_En18
  input [18:0] Wgt_1_362, // sfix19_En18
  input [18:0] Wgt_1_363, // sfix19_En18
  input [18:0] Wgt_1_364, // sfix19_En18
  input [18:0] Wgt_1_365, // sfix19_En18
  input [18:0] Wgt_1_366, // sfix19_En18
  input [18:0] Wgt_1_367, // sfix19_En18
  input [18:0] Wgt_1_368, // sfix19_En18
  input [18:0] Wgt_1_369, // sfix19_En18
  input [18:0] Wgt_1_370, // sfix19_En18
  input [18:0] Wgt_1_371, // sfix19_En18
  input [18:0] Wgt_1_372, // sfix19_En18
  input [18:0] Wgt_1_373, // sfix19_En18
  input [18:0] Wgt_1_374, // sfix19_En18
  input [18:0] Wgt_1_375, // sfix19_En18
  input [18:0] Wgt_1_376, // sfix19_En18
  input [18:0] Wgt_1_377, // sfix19_En18
  input [18:0] Wgt_1_378, // sfix19_En18
  input [18:0] Wgt_1_379, // sfix19_En18
  input [18:0] Wgt_1_380, // sfix19_En18
  input [18:0] Wgt_1_381, // sfix19_En18
  input [18:0] Wgt_1_382, // sfix19_En18
  input [18:0] Wgt_1_383, // sfix19_En18
  input [18:0] Wgt_1_384, // sfix19_En18
  input [18:0] Wgt_1_385, // sfix19_En18
  input [18:0] Wgt_1_386, // sfix19_En18
  input [18:0] Wgt_1_387, // sfix19_En18
  input [18:0] Wgt_1_388, // sfix19_En18
  input [18:0] Wgt_1_389, // sfix19_En18
  input [18:0] Wgt_1_390, // sfix19_En18
  input [18:0] Wgt_1_391, // sfix19_En18
  input [18:0] Wgt_1_392, // sfix19_En18
  input [18:0] Wgt_1_393, // sfix19_En18
  input [18:0] Wgt_1_394, // sfix19_En18
  input [18:0] Wgt_1_395, // sfix19_En18
  input [18:0] Wgt_1_396, // sfix19_En18
  input [18:0] Wgt_1_397, // sfix19_En18
  input [18:0] Wgt_1_398, // sfix19_En18
  input [18:0] Wgt_1_399, // sfix19_En18
  input [18:0] Wgt_1_400, // sfix19_En18
  input [18:0] Wgt_1_401, // sfix19_En18
  input [18:0] Wgt_1_402, // sfix19_En18
  input [18:0] Wgt_1_403, // sfix19_En18
  input [18:0] Wgt_1_404, // sfix19_En18
  input [18:0] Wgt_1_405, // sfix19_En18
  input [18:0] Wgt_1_406, // sfix19_En18
  input [18:0] Wgt_1_407, // sfix19_En18
  input [18:0] Wgt_1_408, // sfix19_En18
  input [18:0] Wgt_1_409, // sfix19_En18
  input [18:0] Wgt_1_410, // sfix19_En18
  input [18:0] Wgt_1_411, // sfix19_En18
  input [18:0] Wgt_1_412, // sfix19_En18
  input [18:0] Wgt_1_413, // sfix19_En18
  input [18:0] Wgt_1_414, // sfix19_En18
  input [18:0] Wgt_1_415, // sfix19_En18
  input [18:0] Wgt_1_416, // sfix19_En18
  input [18:0] Wgt_1_417, // sfix19_En18
  input [18:0] Wgt_1_418, // sfix19_En18
  input [18:0] Wgt_1_419, // sfix19_En18
  input [18:0] Wgt_1_420, // sfix19_En18
  input [18:0] Wgt_1_421, // sfix19_En18
  input [18:0] Wgt_1_422, // sfix19_En18
  input [18:0] Wgt_1_423, // sfix19_En18
  input [18:0] Wgt_1_424, // sfix19_En18
  input [18:0] Wgt_1_425, // sfix19_En18
  input [18:0] Wgt_1_426, // sfix19_En18
  input [18:0] Wgt_1_427, // sfix19_En18
  input [18:0] Wgt_1_428, // sfix19_En18
  input [18:0] Wgt_1_429, // sfix19_En18
  input [18:0] Wgt_1_430, // sfix19_En18
  input [18:0] Wgt_1_431, // sfix19_En18
  input [18:0] Wgt_1_432, // sfix19_En18
  input [18:0] Wgt_1_433, // sfix19_En18
  input [18:0] Wgt_1_434, // sfix19_En18
  input [18:0] Wgt_1_435, // sfix19_En18
  input [18:0] Wgt_1_436, // sfix19_En18
  input [18:0] Wgt_1_437, // sfix19_En18
  input [18:0] Wgt_1_438, // sfix19_En18
  input [18:0] Wgt_1_439, // sfix19_En18
  input [18:0] Wgt_1_440, // sfix19_En18
  input [18:0] Wgt_1_441, // sfix19_En18
  input [18:0] Wgt_1_442, // sfix19_En18
  input [18:0] Wgt_1_443, // sfix19_En18
  input [18:0] Wgt_1_444, // sfix19_En18
  input [18:0] Wgt_1_445, // sfix19_En18
  input [18:0] Wgt_1_446, // sfix19_En18
  input [18:0] Wgt_1_447, // sfix19_En18
  input [18:0] Wgt_1_448, // sfix19_En18
  input [18:0] Wgt_1_449, // sfix19_En18
  input [18:0] Wgt_1_450, // sfix19_En18
  input [18:0] Wgt_1_451, // sfix19_En18
  input [18:0] Wgt_1_452, // sfix19_En18
  input [18:0] Wgt_1_453, // sfix19_En18
  input [18:0] Wgt_1_454, // sfix19_En18
  input [18:0] Wgt_1_455, // sfix19_En18
  input [18:0] Wgt_1_456, // sfix19_En18
  input [18:0] Wgt_1_457, // sfix19_En18
  input [18:0] Wgt_1_458, // sfix19_En18
  input [18:0] Wgt_1_459, // sfix19_En18
  input [18:0] Wgt_1_460, // sfix19_En18
  input [18:0] Wgt_1_461, // sfix19_En18
  input [18:0] Wgt_1_462, // sfix19_En18
  input [18:0] Wgt_1_463, // sfix19_En18
  input [18:0] Wgt_1_464, // sfix19_En18
  input [18:0] Wgt_1_465, // sfix19_En18
  input [18:0] Wgt_1_466, // sfix19_En18
  input [18:0] Wgt_1_467, // sfix19_En18
  input [18:0] Wgt_1_468, // sfix19_En18
  input [18:0] Wgt_1_469, // sfix19_En18
  input [18:0] Wgt_1_470, // sfix19_En18
  input [18:0] Wgt_1_471, // sfix19_En18
  input [18:0] Wgt_1_472, // sfix19_En18
  input [18:0] Wgt_1_473, // sfix19_En18
  input [18:0] Wgt_1_474, // sfix19_En18
  input [18:0] Wgt_1_475, // sfix19_En18
  input [18:0] Wgt_1_476, // sfix19_En18
  input [18:0] Wgt_1_477, // sfix19_En18
  input [18:0] Wgt_1_478, // sfix19_En18
  input [18:0] Wgt_1_479, // sfix19_En18
  input [18:0] Wgt_1_480, // sfix19_En18
  input [18:0] Wgt_1_481, // sfix19_En18
  input [18:0] Wgt_1_482, // sfix19_En18
  input [18:0] Wgt_1_483, // sfix19_En18
  input [18:0] Wgt_1_484, // sfix19_En18
  input [18:0] Wgt_1_485, // sfix19_En18
  input [18:0] Wgt_1_486, // sfix19_En18
  input [18:0] Wgt_1_487, // sfix19_En18
  input [18:0] Wgt_1_488, // sfix19_En18
  input [18:0] Wgt_1_489, // sfix19_En18
  input [18:0] Wgt_1_490, // sfix19_En18
  input [18:0] Wgt_1_491, // sfix19_En18
  input [18:0] Wgt_1_492, // sfix19_En18
  input [18:0] Wgt_1_493, // sfix19_En18
  input [18:0] Wgt_1_494, // sfix19_En18
  input [18:0] Wgt_1_495, // sfix19_En18
  input [18:0] Wgt_1_496, // sfix19_En18
  input [18:0] Wgt_1_497, // sfix19_En18
  input [18:0] Wgt_1_498, // sfix19_En18
  input [18:0] Wgt_1_499, // sfix19_En18
  input [18:0] Wgt_1_500, // sfix19_En18
  input [18:0] Wgt_1_501, // sfix19_En18
  input [18:0] Wgt_1_502, // sfix19_En18
  input [18:0] Wgt_1_503, // sfix19_En18
  input [18:0] Wgt_1_504, // sfix19_En18
  input [18:0] Wgt_1_505, // sfix19_En18
  input [18:0] Wgt_1_506, // sfix19_En18
  input [18:0] Wgt_1_507, // sfix19_En18
  input [18:0] Wgt_1_508, // sfix19_En18
  input [18:0] Wgt_1_509, // sfix19_En18
  input [18:0] Wgt_1_510, // sfix19_En18
  input [18:0] Wgt_1_511, // sfix19_En18
  input [18:0] Wgt_1_512, // sfix19_En18
  input [18:0] Wgt_1_513, // sfix19_En18
  input [18:0] Wgt_1_514, // sfix19_En18
  input [18:0] Wgt_1_515, // sfix19_En18
  input [18:0] Wgt_1_516, // sfix19_En18
  input [18:0] Wgt_1_517, // sfix19_En18
  input [18:0] Wgt_1_518, // sfix19_En18
  input [18:0] Wgt_1_519, // sfix19_En18
  input [18:0] Wgt_1_520, // sfix19_En18
  input [18:0] Wgt_1_521, // sfix19_En18
  input [18:0] Wgt_1_522, // sfix19_En18
  input [18:0] Wgt_1_523, // sfix19_En18
  input [18:0] Wgt_1_524, // sfix19_En18
  input [18:0] Wgt_1_525, // sfix19_En18
  input [18:0] Wgt_1_526, // sfix19_En18
  input [18:0] Wgt_1_527, // sfix19_En18
  input [18:0] Wgt_1_528, // sfix19_En18
  input [18:0] Wgt_1_529, // sfix19_En18
  input [18:0] Wgt_1_530, // sfix19_En18
  input [18:0] Wgt_1_531, // sfix19_En18
  input [18:0] Wgt_1_532, // sfix19_En18
  input [18:0] Wgt_1_533, // sfix19_En18
  input [18:0] Wgt_1_534, // sfix19_En18
  input [18:0] Wgt_1_535, // sfix19_En18
  input [18:0] Wgt_1_536, // sfix19_En18
  input [18:0] Wgt_1_537, // sfix19_En18
  input [18:0] Wgt_1_538, // sfix19_En18
  input [18:0] Wgt_1_539, // sfix19_En18
  input [18:0] Wgt_1_540, // sfix19_En18
  input [18:0] Wgt_1_541, // sfix19_En18
  input [18:0] Wgt_1_542, // sfix19_En18
  input [18:0] Wgt_1_543, // sfix19_En18
  input [18:0] Wgt_1_544, // sfix19_En18
  input [18:0] Wgt_1_545, // sfix19_En18
  input [18:0] Wgt_1_546, // sfix19_En18
  input [18:0] Wgt_1_547, // sfix19_En18
  input [18:0] Wgt_1_548, // sfix19_En18
  input [18:0] Wgt_1_549, // sfix19_En18
  input [18:0] Wgt_1_550, // sfix19_En18
  input [18:0] Wgt_1_551, // sfix19_En18
  input [18:0] Wgt_1_552, // sfix19_En18
  input [18:0] Wgt_1_553, // sfix19_En18
  input [18:0] Wgt_1_554, // sfix19_En18
  input [18:0] Wgt_1_555, // sfix19_En18
  input [18:0] Wgt_1_556, // sfix19_En18
  input [18:0] Wgt_1_557, // sfix19_En18
  input [18:0] Wgt_1_558, // sfix19_En18
  input [18:0] Wgt_1_559, // sfix19_En18
  input [18:0] Wgt_1_560, // sfix19_En18
  input [18:0] Wgt_1_561, // sfix19_En18
  input [18:0] Wgt_1_562, // sfix19_En18
  input [18:0] Wgt_1_563, // sfix19_En18
  input [18:0] Wgt_1_564, // sfix19_En18
  input [18:0] Wgt_1_565, // sfix19_En18
  input [18:0] Wgt_1_566, // sfix19_En18
  input [18:0] Wgt_1_567, // sfix19_En18
  input [18:0] Wgt_1_568, // sfix19_En18
  input [18:0] Wgt_1_569, // sfix19_En18
  input [18:0] Wgt_1_570, // sfix19_En18
  input [18:0] Wgt_1_571, // sfix19_En18
  input [18:0] Wgt_1_572, // sfix19_En18
  input [18:0] Wgt_1_573, // sfix19_En18
  input [18:0] Wgt_1_574, // sfix19_En18
  input [18:0] Wgt_1_575, // sfix19_En18
  input [18:0] Wgt_1_576, // sfix19_En18
  input [18:0] Wgt_1_577, // sfix19_En18
  input [18:0] Wgt_1_578, // sfix19_En18
  input [18:0] Wgt_1_579, // sfix19_En18
  input [18:0] Wgt_1_580, // sfix19_En18
  input [18:0] Wgt_1_581, // sfix19_En18
  input [18:0] Wgt_1_582, // sfix19_En18
  input [18:0] Wgt_1_583, // sfix19_En18
  input [18:0] Wgt_1_584, // sfix19_En18
  input [18:0] Wgt_1_585, // sfix19_En18
  input [18:0] Wgt_1_586, // sfix19_En18
  input [18:0] Wgt_1_587, // sfix19_En18
  input [18:0] Wgt_1_588, // sfix19_En18
  input [18:0] Wgt_1_589, // sfix19_En18
  input [18:0] Wgt_1_590, // sfix19_En18
  input [18:0] Wgt_1_591, // sfix19_En18
  input [18:0] Wgt_1_592, // sfix19_En18
  input [18:0] Wgt_1_593, // sfix19_En18
  input [18:0] Wgt_1_594, // sfix19_En18
  input [18:0] Wgt_1_595, // sfix19_En18
  input [18:0] Wgt_1_596, // sfix19_En18
  input [18:0] Wgt_1_597, // sfix19_En18
  input [18:0] Wgt_1_598, // sfix19_En18
  input [18:0] Wgt_1_599, // sfix19_En18
  input [18:0] Wgt_1_600, // sfix19_En18
  input [18:0] Wgt_1_601, // sfix19_En18
  input [18:0] Wgt_1_602, // sfix19_En18
  input [18:0] Wgt_1_603, // sfix19_En18
  input [18:0] Wgt_1_604, // sfix19_En18
  input [18:0] Wgt_1_605, // sfix19_En18
  input [18:0] Wgt_1_606, // sfix19_En18
  input [18:0] Wgt_1_607, // sfix19_En18
  input [18:0] Wgt_1_608, // sfix19_En18
  input [18:0] Wgt_1_609, // sfix19_En18
  input [18:0] Wgt_1_610, // sfix19_En18
  input [18:0] Wgt_1_611, // sfix19_En18
  input [18:0] Wgt_1_612, // sfix19_En18
  input [18:0] Wgt_1_613, // sfix19_En18
  input [18:0] Wgt_1_614, // sfix19_En18
  input [18:0] Wgt_1_615, // sfix19_En18
  input [18:0] Wgt_1_616, // sfix19_En18
  input [18:0] Wgt_1_617, // sfix19_En18
  input [18:0] Wgt_1_618, // sfix19_En18
  input [18:0] Wgt_1_619, // sfix19_En18
  input [18:0] Wgt_1_620, // sfix19_En18
  input [18:0] Wgt_1_621, // sfix19_En18
  input [18:0] Wgt_1_622, // sfix19_En18
  input [18:0] Wgt_1_623, // sfix19_En18
  input [18:0] Wgt_1_624, // sfix19_En18
  input [18:0] Wgt_1_625, // sfix19_En18
  input [18:0] Wgt_1_626, // sfix19_En18
  input [18:0] Wgt_1_627, // sfix19_En18
  input [18:0] Wgt_1_628, // sfix19_En18
  input [18:0] Wgt_1_629, // sfix19_En18
  input [18:0] Wgt_1_630, // sfix19_En18
  input [18:0] Wgt_1_631, // sfix19_En18
  input [18:0] Wgt_1_632, // sfix19_En18
  input [18:0] Wgt_1_633, // sfix19_En18
  input [18:0] Wgt_1_634, // sfix19_En18
  input [18:0] Wgt_1_635, // sfix19_En18
  input [18:0] Wgt_1_636, // sfix19_En18
  input [18:0] Wgt_1_637, // sfix19_En18
  input [18:0] Wgt_1_638, // sfix19_En18
  input [18:0] Wgt_1_639, // sfix19_En18
  input [18:0] Wgt_1_640, // sfix19_En18
  input [18:0] Wgt_1_641, // sfix19_En18
  input [18:0] Wgt_1_642, // sfix19_En18
  input [18:0] Wgt_1_643, // sfix19_En18
  input [18:0] Wgt_1_644, // sfix19_En18
  input [18:0] Wgt_1_645, // sfix19_En18
  input [18:0] Wgt_1_646, // sfix19_En18
  input [18:0] Wgt_1_647, // sfix19_En18
  input [18:0] Wgt_1_648, // sfix19_En18
  input [18:0] Wgt_1_649, // sfix19_En18
  input [18:0] Wgt_1_650, // sfix19_En18
  input [18:0] Wgt_1_651, // sfix19_En18
  input [18:0] Wgt_1_652, // sfix19_En18
  input [18:0] Wgt_1_653, // sfix19_En18
  input [18:0] Wgt_1_654, // sfix19_En18
  input [18:0] Wgt_1_655, // sfix19_En18
  input [18:0] Wgt_1_656, // sfix19_En18
  input [18:0] Wgt_1_657, // sfix19_En18
  input [18:0] Wgt_1_658, // sfix19_En18
  input [18:0] Wgt_1_659, // sfix19_En18
  input [18:0] Wgt_1_660, // sfix19_En18
  input [18:0] Wgt_1_661, // sfix19_En18
  input [18:0] Wgt_1_662, // sfix19_En18
  input [18:0] Wgt_1_663, // sfix19_En18
  input [18:0] Wgt_1_664, // sfix19_En18
  input [18:0] Wgt_1_665, // sfix19_En18
  input [18:0] Wgt_1_666, // sfix19_En18
  input [18:0] Wgt_1_667, // sfix19_En18
  input [18:0] Wgt_1_668, // sfix19_En18
  input [18:0] Wgt_1_669, // sfix19_En18
  input [18:0] Wgt_1_670, // sfix19_En18
  input [18:0] Wgt_1_671, // sfix19_En18
  input [18:0] Wgt_1_672, // sfix19_En18
  input [18:0] Wgt_1_673, // sfix19_En18
  input [18:0] Wgt_1_674, // sfix19_En18
  input [18:0] Wgt_1_675, // sfix19_En18
  input [18:0] Wgt_1_676, // sfix19_En18
  input [18:0] Wgt_1_677, // sfix19_En18
  input [18:0] Wgt_1_678, // sfix19_En18
  input [18:0] Wgt_1_679, // sfix19_En18
  input [18:0] Wgt_1_680, // sfix19_En18
  input [18:0] Wgt_1_681, // sfix19_En18
  input [18:0] Wgt_1_682, // sfix19_En18
  input [18:0] Wgt_1_683, // sfix19_En18
  input [18:0] Wgt_1_684, // sfix19_En18
  input [18:0] Wgt_1_685, // sfix19_En18
  input [18:0] Wgt_1_686, // sfix19_En18
  input [18:0] Wgt_1_687, // sfix19_En18
  input [18:0] Wgt_1_688, // sfix19_En18
  input [18:0] Wgt_1_689, // sfix19_En18
  input [18:0] Wgt_1_690, // sfix19_En18
  input [18:0] Wgt_1_691, // sfix19_En18
  input [18:0] Wgt_1_692, // sfix19_En18
  input [18:0] Wgt_1_693, // sfix19_En18
  input [18:0] Wgt_1_694, // sfix19_En18
  input [18:0] Wgt_1_695, // sfix19_En18
  input [18:0] Wgt_1_696, // sfix19_En18
  input [18:0] Wgt_1_697, // sfix19_En18
  input [18:0] Wgt_1_698, // sfix19_En18
  input [18:0] Wgt_1_699, // sfix19_En18
  input [18:0] Wgt_1_700, // sfix19_En18
  input [18:0] Wgt_1_701, // sfix19_En18
  input [18:0] Wgt_1_702, // sfix19_En18
  input [18:0] Wgt_1_703, // sfix19_En18
  input [18:0] Wgt_1_704, // sfix19_En18
  input [18:0] Wgt_1_705, // sfix19_En18
  input [18:0] Wgt_1_706, // sfix19_En18
  input [18:0] Wgt_1_707, // sfix19_En18
  input [18:0] Wgt_1_708, // sfix19_En18
  input [18:0] Wgt_1_709, // sfix19_En18
  input [18:0] Wgt_1_710, // sfix19_En18
  input [18:0] Wgt_1_711, // sfix19_En18
  input [18:0] Wgt_1_712, // sfix19_En18
  input [18:0] Wgt_1_713, // sfix19_En18
  input [18:0] Wgt_1_714, // sfix19_En18
  input [18:0] Wgt_1_715, // sfix19_En18
  input [18:0] Wgt_1_716, // sfix19_En18
  input [18:0] Wgt_1_717, // sfix19_En18
  input [18:0] Wgt_1_718, // sfix19_En18
  input [18:0] Wgt_1_719, // sfix19_En18
  input [18:0] Wgt_1_720, // sfix19_En18
  input [18:0] Wgt_1_721, // sfix19_En18
  input [18:0] Wgt_1_722, // sfix19_En18
  input [18:0] Wgt_1_723, // sfix19_En18
  input [18:0] Wgt_1_724, // sfix19_En18
  input [18:0] Wgt_1_725, // sfix19_En18
  input [18:0] Wgt_1_726, // sfix19_En18
  input [18:0] Wgt_1_727, // sfix19_En18
  input [18:0] Wgt_1_728, // sfix19_En18
  input [18:0] Wgt_1_729, // sfix19_En18
  input [18:0] Wgt_1_730, // sfix19_En18
  input [18:0] Wgt_1_731, // sfix19_En18
  input [18:0] Wgt_1_732, // sfix19_En18
  input [18:0] Wgt_1_733, // sfix19_En18
  input [18:0] Wgt_1_734, // sfix19_En18
  input [18:0] Wgt_1_735, // sfix19_En18
  input [18:0] Wgt_1_736, // sfix19_En18
  input [18:0] Wgt_1_737, // sfix19_En18
  input [18:0] Wgt_1_738, // sfix19_En18
  input [18:0] Wgt_1_739, // sfix19_En18
  input [18:0] Wgt_1_740, // sfix19_En18
  input [18:0] Wgt_1_741, // sfix19_En18
  input [18:0] Wgt_1_742, // sfix19_En18
  input [18:0] Wgt_1_743, // sfix19_En18
  input [18:0] Wgt_1_744, // sfix19_En18
  input [18:0] Wgt_1_745, // sfix19_En18
  input [18:0] Wgt_1_746, // sfix19_En18
  input [18:0] Wgt_1_747, // sfix19_En18
  input [18:0] Wgt_1_748, // sfix19_En18
  input [18:0] Wgt_1_749, // sfix19_En18
  input [18:0] Wgt_1_750, // sfix19_En18
  input [18:0] Wgt_1_751, // sfix19_En18
  input [18:0] Wgt_1_752, // sfix19_En18
  input [18:0] Wgt_1_753, // sfix19_En18
  input [18:0] Wgt_1_754, // sfix19_En18
  input [18:0] Wgt_1_755, // sfix19_En18
  input [18:0] Wgt_1_756, // sfix19_En18
  input [18:0] Wgt_1_757, // sfix19_En18
  input [18:0] Wgt_1_758, // sfix19_En18
  input [18:0] Wgt_1_759, // sfix19_En18
  input [18:0] Wgt_1_760, // sfix19_En18
  input [18:0] Wgt_1_761, // sfix19_En18
  input [18:0] Wgt_1_762, // sfix19_En18
  input [18:0] Wgt_1_763, // sfix19_En18
  input [18:0] Wgt_1_764, // sfix19_En18
  input [18:0] Wgt_1_765, // sfix19_En18
  input [18:0] Wgt_1_766, // sfix19_En18
  input [18:0] Wgt_1_767, // sfix19_En18
  input [18:0] Wgt_1_768, // sfix19_En18
  input [18:0] Wgt_1_769, // sfix19_En18
  input [18:0] Wgt_1_770, // sfix19_En18
  input [18:0] Wgt_1_771, // sfix19_En18
  input [18:0] Wgt_1_772, // sfix19_En18
  input [18:0] Wgt_1_773, // sfix19_En18
  input [18:0] Wgt_1_774, // sfix19_En18
  input [18:0] Wgt_1_775, // sfix19_En18
  input [18:0] Wgt_1_776, // sfix19_En18
  input [18:0] Wgt_1_777, // sfix19_En18
  input [18:0] Wgt_1_778, // sfix19_En18
  input [18:0] Wgt_1_779, // sfix19_En18
  input [18:0] Wgt_1_780, // sfix19_En18
  input [18:0] Wgt_1_781, // sfix19_En18
  input [18:0] Wgt_1_782, // sfix19_En18
  input [18:0] Wgt_1_783, // sfix19_En18
  input [18:0] Wgt_1_784, // sfix19_En18
  input [18:0] Wgt_2_0, // sfix19_En18
  input [18:0] Wgt_2_1, // sfix19_En18
  input [18:0] Wgt_2_2, // sfix19_En18
  input [18:0] Wgt_2_3, // sfix19_En18
  input [18:0] Wgt_2_4, // sfix19_En18
  input [18:0] Wgt_2_5, // sfix19_En18
  input [18:0] Wgt_2_6, // sfix19_En18
  input [18:0] Wgt_2_7, // sfix19_En18
  input [18:0] Wgt_2_8, // sfix19_En18
  input [18:0] Wgt_2_9, // sfix19_En18
  input [18:0] Wgt_2_10, // sfix19_En18
  input [18:0] Wgt_2_11, // sfix19_En18
  input [18:0] Wgt_2_12, // sfix19_En18
  input [18:0] Wgt_2_13, // sfix19_En18
  input [18:0] Wgt_2_14, // sfix19_En18
  input [18:0] Wgt_2_15, // sfix19_En18
  input [18:0] Wgt_2_16, // sfix19_En18
  input [18:0] Wgt_2_17, // sfix19_En18
  input [18:0] Wgt_2_18, // sfix19_En18
  input [18:0] Wgt_2_19, // sfix19_En18
  input [18:0] Wgt_2_20, // sfix19_En18
  input [18:0] Wgt_2_21, // sfix19_En18
  input [18:0] Wgt_2_22, // sfix19_En18
  input [18:0] Wgt_2_23, // sfix19_En18
  input [18:0] Wgt_2_24, // sfix19_En18
  input [18:0] Wgt_2_25, // sfix19_En18
  input [18:0] Wgt_2_26, // sfix19_En18
  input [18:0] Wgt_2_27, // sfix19_En18
  input [18:0] Wgt_2_28, // sfix19_En18
  input [18:0] Wgt_2_29, // sfix19_En18
  input [18:0] Wgt_2_30, // sfix19_En18
  input [18:0] Wgt_2_31, // sfix19_En18
  input [18:0] Wgt_2_32, // sfix19_En18
  input [18:0] Wgt_2_33, // sfix19_En18
  input [18:0] Wgt_2_34, // sfix19_En18
  input [18:0] Wgt_2_35, // sfix19_En18
  input [18:0] Wgt_2_36, // sfix19_En18
  input [18:0] Wgt_2_37, // sfix19_En18
  input [18:0] Wgt_2_38, // sfix19_En18
  input [18:0] Wgt_2_39, // sfix19_En18
  input [18:0] Wgt_2_40, // sfix19_En18
  input [18:0] Wgt_2_41, // sfix19_En18
  input [18:0] Wgt_2_42, // sfix19_En18
  input [18:0] Wgt_2_43, // sfix19_En18
  input [18:0] Wgt_2_44, // sfix19_En18
  input [18:0] Wgt_2_45, // sfix19_En18
  input [18:0] Wgt_2_46, // sfix19_En18
  input [18:0] Wgt_2_47, // sfix19_En18
  input [18:0] Wgt_2_48, // sfix19_En18
  input [18:0] Wgt_2_49, // sfix19_En18
  input [18:0] Wgt_2_50, // sfix19_En18
  input [18:0] Wgt_2_51, // sfix19_En18
  input [18:0] Wgt_2_52, // sfix19_En18
  input [18:0] Wgt_2_53, // sfix19_En18
  input [18:0] Wgt_2_54, // sfix19_En18
  input [18:0] Wgt_2_55, // sfix19_En18
  input [18:0] Wgt_2_56, // sfix19_En18
  input [18:0] Wgt_2_57, // sfix19_En18
  input [18:0] Wgt_2_58, // sfix19_En18
  input [18:0] Wgt_2_59, // sfix19_En18
  input [18:0] Wgt_2_60, // sfix19_En18
  input [18:0] Wgt_2_61, // sfix19_En18
  input [18:0] Wgt_2_62, // sfix19_En18
  input [18:0] Wgt_2_63, // sfix19_En18
  input [18:0] Wgt_2_64, // sfix19_En18
  input [18:0] Wgt_2_65, // sfix19_En18
  input [18:0] Wgt_2_66, // sfix19_En18
  input [18:0] Wgt_2_67, // sfix19_En18
  input [18:0] Wgt_2_68, // sfix19_En18
  input [18:0] Wgt_2_69, // sfix19_En18
  input [18:0] Wgt_2_70, // sfix19_En18
  input [18:0] Wgt_2_71, // sfix19_En18
  input [18:0] Wgt_2_72, // sfix19_En18
  input [18:0] Wgt_2_73, // sfix19_En18
  input [18:0] Wgt_2_74, // sfix19_En18
  input [18:0] Wgt_2_75, // sfix19_En18
  input [18:0] Wgt_2_76, // sfix19_En18
  input [18:0] Wgt_2_77, // sfix19_En18
  input [18:0] Wgt_2_78, // sfix19_En18
  input [18:0] Wgt_2_79, // sfix19_En18
  input [18:0] Wgt_2_80, // sfix19_En18
  input [18:0] Wgt_2_81, // sfix19_En18
  input [18:0] Wgt_2_82, // sfix19_En18
  input [18:0] Wgt_2_83, // sfix19_En18
  input [18:0] Wgt_2_84, // sfix19_En18
  input [18:0] Wgt_2_85, // sfix19_En18
  input [18:0] Wgt_2_86, // sfix19_En18
  input [18:0] Wgt_2_87, // sfix19_En18
  input [18:0] Wgt_2_88, // sfix19_En18
  input [18:0] Wgt_2_89, // sfix19_En18
  input [18:0] Wgt_2_90, // sfix19_En18
  input [18:0] Wgt_2_91, // sfix19_En18
  input [18:0] Wgt_2_92, // sfix19_En18
  input [18:0] Wgt_2_93, // sfix19_En18
  input [18:0] Wgt_2_94, // sfix19_En18
  input [18:0] Wgt_2_95, // sfix19_En18
  input [18:0] Wgt_2_96, // sfix19_En18
  input [18:0] Wgt_2_97, // sfix19_En18
  input [18:0] Wgt_2_98, // sfix19_En18
  input [18:0] Wgt_2_99, // sfix19_En18
  input [18:0] Wgt_2_100, // sfix19_En18
  input [18:0] Wgt_2_101, // sfix19_En18
  input [18:0] Wgt_2_102, // sfix19_En18
  input [18:0] Wgt_2_103, // sfix19_En18
  input [18:0] Wgt_2_104, // sfix19_En18
  input [18:0] Wgt_2_105, // sfix19_En18
  input [18:0] Wgt_2_106, // sfix19_En18
  input [18:0] Wgt_2_107, // sfix19_En18
  input [18:0] Wgt_2_108, // sfix19_En18
  input [18:0] Wgt_2_109, // sfix19_En18
  input [18:0] Wgt_2_110, // sfix19_En18
  input [18:0] Wgt_2_111, // sfix19_En18
  input [18:0] Wgt_2_112, // sfix19_En18
  input [18:0] Wgt_2_113, // sfix19_En18
  input [18:0] Wgt_2_114, // sfix19_En18
  input [18:0] Wgt_2_115, // sfix19_En18
  input [18:0] Wgt_2_116, // sfix19_En18
  input [18:0] Wgt_2_117, // sfix19_En18
  input [18:0] Wgt_2_118, // sfix19_En18
  input [18:0] Wgt_2_119, // sfix19_En18
  input [18:0] Wgt_2_120, // sfix19_En18
  input [18:0] Wgt_2_121, // sfix19_En18
  input [18:0] Wgt_2_122, // sfix19_En18
  input [18:0] Wgt_2_123, // sfix19_En18
  input [18:0] Wgt_2_124, // sfix19_En18
  input [18:0] Wgt_2_125, // sfix19_En18
  input [18:0] Wgt_2_126, // sfix19_En18
  input [18:0] Wgt_2_127, // sfix19_En18
  input [18:0] Wgt_2_128, // sfix19_En18
  input [18:0] Wgt_2_129, // sfix19_En18
  input [18:0] Wgt_2_130, // sfix19_En18
  input [18:0] Wgt_2_131, // sfix19_En18
  input [18:0] Wgt_2_132, // sfix19_En18
  input [18:0] Wgt_2_133, // sfix19_En18
  input [18:0] Wgt_2_134, // sfix19_En18
  input [18:0] Wgt_2_135, // sfix19_En18
  input [18:0] Wgt_2_136, // sfix19_En18
  input [18:0] Wgt_2_137, // sfix19_En18
  input [18:0] Wgt_2_138, // sfix19_En18
  input [18:0] Wgt_2_139, // sfix19_En18
  input [18:0] Wgt_2_140, // sfix19_En18
  input [18:0] Wgt_2_141, // sfix19_En18
  input [18:0] Wgt_2_142, // sfix19_En18
  input [18:0] Wgt_2_143, // sfix19_En18
  input [18:0] Wgt_2_144, // sfix19_En18
  input [18:0] Wgt_2_145, // sfix19_En18
  input [18:0] Wgt_2_146, // sfix19_En18
  input [18:0] Wgt_2_147, // sfix19_En18
  input [18:0] Wgt_2_148, // sfix19_En18
  input [18:0] Wgt_2_149, // sfix19_En18
  input [18:0] Wgt_2_150, // sfix19_En18
  input [18:0] Wgt_2_151, // sfix19_En18
  input [18:0] Wgt_2_152, // sfix19_En18
  input [18:0] Wgt_2_153, // sfix19_En18
  input [18:0] Wgt_2_154, // sfix19_En18
  input [18:0] Wgt_2_155, // sfix19_En18
  input [18:0] Wgt_2_156, // sfix19_En18
  input [18:0] Wgt_2_157, // sfix19_En18
  input [18:0] Wgt_2_158, // sfix19_En18
  input [18:0] Wgt_2_159, // sfix19_En18
  input [18:0] Wgt_2_160, // sfix19_En18
  input [18:0] Wgt_2_161, // sfix19_En18
  input [18:0] Wgt_2_162, // sfix19_En18
  input [18:0] Wgt_2_163, // sfix19_En18
  input [18:0] Wgt_2_164, // sfix19_En18
  input [18:0] Wgt_2_165, // sfix19_En18
  input [18:0] Wgt_2_166, // sfix19_En18
  input [18:0] Wgt_2_167, // sfix19_En18
  input [18:0] Wgt_2_168, // sfix19_En18
  input [18:0] Wgt_2_169, // sfix19_En18
  input [18:0] Wgt_2_170, // sfix19_En18
  input [18:0] Wgt_2_171, // sfix19_En18
  input [18:0] Wgt_2_172, // sfix19_En18
  input [18:0] Wgt_2_173, // sfix19_En18
  input [18:0] Wgt_2_174, // sfix19_En18
  input [18:0] Wgt_2_175, // sfix19_En18
  input [18:0] Wgt_2_176, // sfix19_En18
  input [18:0] Wgt_2_177, // sfix19_En18
  input [18:0] Wgt_2_178, // sfix19_En18
  input [18:0] Wgt_2_179, // sfix19_En18
  input [18:0] Wgt_2_180, // sfix19_En18
  input [18:0] Wgt_2_181, // sfix19_En18
  input [18:0] Wgt_2_182, // sfix19_En18
  input [18:0] Wgt_2_183, // sfix19_En18
  input [18:0] Wgt_2_184, // sfix19_En18
  input [18:0] Wgt_2_185, // sfix19_En18
  input [18:0] Wgt_2_186, // sfix19_En18
  input [18:0] Wgt_2_187, // sfix19_En18
  input [18:0] Wgt_2_188, // sfix19_En18
  input [18:0] Wgt_2_189, // sfix19_En18
  input [18:0] Wgt_2_190, // sfix19_En18
  input [18:0] Wgt_2_191, // sfix19_En18
  input [18:0] Wgt_2_192, // sfix19_En18
  input [18:0] Wgt_2_193, // sfix19_En18
  input [18:0] Wgt_2_194, // sfix19_En18
  input [18:0] Wgt_2_195, // sfix19_En18
  input [18:0] Wgt_2_196, // sfix19_En18
  input [18:0] Wgt_2_197, // sfix19_En18
  input [18:0] Wgt_2_198, // sfix19_En18
  input [18:0] Wgt_2_199, // sfix19_En18
  input [18:0] Wgt_2_200, // sfix19_En18
  input [18:0] Wgt_2_201, // sfix19_En18
  input [18:0] Wgt_2_202, // sfix19_En18
  input [18:0] Wgt_2_203, // sfix19_En18
  input [18:0] Wgt_2_204, // sfix19_En18
  input [18:0] Wgt_2_205, // sfix19_En18
  input [18:0] Wgt_2_206, // sfix19_En18
  input [18:0] Wgt_2_207, // sfix19_En18
  input [18:0] Wgt_2_208, // sfix19_En18
  input [18:0] Wgt_2_209, // sfix19_En18
  input [18:0] Wgt_2_210, // sfix19_En18
  input [18:0] Wgt_2_211, // sfix19_En18
  input [18:0] Wgt_2_212, // sfix19_En18
  input [18:0] Wgt_2_213, // sfix19_En18
  input [18:0] Wgt_2_214, // sfix19_En18
  input [18:0] Wgt_2_215, // sfix19_En18
  input [18:0] Wgt_2_216, // sfix19_En18
  input [18:0] Wgt_2_217, // sfix19_En18
  input [18:0] Wgt_2_218, // sfix19_En18
  input [18:0] Wgt_2_219, // sfix19_En18
  input [18:0] Wgt_2_220, // sfix19_En18
  input [18:0] Wgt_2_221, // sfix19_En18
  input [18:0] Wgt_2_222, // sfix19_En18
  input [18:0] Wgt_2_223, // sfix19_En18
  input [18:0] Wgt_2_224, // sfix19_En18
  input [18:0] Wgt_2_225, // sfix19_En18
  input [18:0] Wgt_2_226, // sfix19_En18
  input [18:0] Wgt_2_227, // sfix19_En18
  input [18:0] Wgt_2_228, // sfix19_En18
  input [18:0] Wgt_2_229, // sfix19_En18
  input [18:0] Wgt_2_230, // sfix19_En18
  input [18:0] Wgt_2_231, // sfix19_En18
  input [18:0] Wgt_2_232, // sfix19_En18
  input [18:0] Wgt_2_233, // sfix19_En18
  input [18:0] Wgt_2_234, // sfix19_En18
  input [18:0] Wgt_2_235, // sfix19_En18
  input [18:0] Wgt_2_236, // sfix19_En18
  input [18:0] Wgt_2_237, // sfix19_En18
  input [18:0] Wgt_2_238, // sfix19_En18
  input [18:0] Wgt_2_239, // sfix19_En18
  input [18:0] Wgt_2_240, // sfix19_En18
  input [18:0] Wgt_2_241, // sfix19_En18
  input [18:0] Wgt_2_242, // sfix19_En18
  input [18:0] Wgt_2_243, // sfix19_En18
  input [18:0] Wgt_2_244, // sfix19_En18
  input [18:0] Wgt_2_245, // sfix19_En18
  input [18:0] Wgt_2_246, // sfix19_En18
  input [18:0] Wgt_2_247, // sfix19_En18
  input [18:0] Wgt_2_248, // sfix19_En18
  input [18:0] Wgt_2_249, // sfix19_En18
  input [18:0] Wgt_2_250, // sfix19_En18
  input [18:0] Wgt_2_251, // sfix19_En18
  input [18:0] Wgt_2_252, // sfix19_En18
  input [18:0] Wgt_2_253, // sfix19_En18
  input [18:0] Wgt_2_254, // sfix19_En18
  input [18:0] Wgt_2_255, // sfix19_En18
  input [18:0] Wgt_2_256, // sfix19_En18
  input [18:0] Wgt_2_257, // sfix19_En18
  input [18:0] Wgt_2_258, // sfix19_En18
  input [18:0] Wgt_2_259, // sfix19_En18
  input [18:0] Wgt_2_260, // sfix19_En18
  input [18:0] Wgt_2_261, // sfix19_En18
  input [18:0] Wgt_2_262, // sfix19_En18
  input [18:0] Wgt_2_263, // sfix19_En18
  input [18:0] Wgt_2_264, // sfix19_En18
  input [18:0] Wgt_2_265, // sfix19_En18
  input [18:0] Wgt_2_266, // sfix19_En18
  input [18:0] Wgt_2_267, // sfix19_En18
  input [18:0] Wgt_2_268, // sfix19_En18
  input [18:0] Wgt_2_269, // sfix19_En18
  input [18:0] Wgt_2_270, // sfix19_En18
  input [18:0] Wgt_2_271, // sfix19_En18
  input [18:0] Wgt_2_272, // sfix19_En18
  input [18:0] Wgt_2_273, // sfix19_En18
  input [18:0] Wgt_2_274, // sfix19_En18
  input [18:0] Wgt_2_275, // sfix19_En18
  input [18:0] Wgt_2_276, // sfix19_En18
  input [18:0] Wgt_2_277, // sfix19_En18
  input [18:0] Wgt_2_278, // sfix19_En18
  input [18:0] Wgt_2_279, // sfix19_En18
  input [18:0] Wgt_2_280, // sfix19_En18
  input [18:0] Wgt_2_281, // sfix19_En18
  input [18:0] Wgt_2_282, // sfix19_En18
  input [18:0] Wgt_2_283, // sfix19_En18
  input [18:0] Wgt_2_284, // sfix19_En18
  input [18:0] Wgt_2_285, // sfix19_En18
  input [18:0] Wgt_2_286, // sfix19_En18
  input [18:0] Wgt_2_287, // sfix19_En18
  input [18:0] Wgt_2_288, // sfix19_En18
  input [18:0] Wgt_2_289, // sfix19_En18
  input [18:0] Wgt_2_290, // sfix19_En18
  input [18:0] Wgt_2_291, // sfix19_En18
  input [18:0] Wgt_2_292, // sfix19_En18
  input [18:0] Wgt_2_293, // sfix19_En18
  input [18:0] Wgt_2_294, // sfix19_En18
  input [18:0] Wgt_2_295, // sfix19_En18
  input [18:0] Wgt_2_296, // sfix19_En18
  input [18:0] Wgt_2_297, // sfix19_En18
  input [18:0] Wgt_2_298, // sfix19_En18
  input [18:0] Wgt_2_299, // sfix19_En18
  input [18:0] Wgt_2_300, // sfix19_En18
  input [18:0] Wgt_2_301, // sfix19_En18
  input [18:0] Wgt_2_302, // sfix19_En18
  input [18:0] Wgt_2_303, // sfix19_En18
  input [18:0] Wgt_2_304, // sfix19_En18
  input [18:0] Wgt_2_305, // sfix19_En18
  input [18:0] Wgt_2_306, // sfix19_En18
  input [18:0] Wgt_2_307, // sfix19_En18
  input [18:0] Wgt_2_308, // sfix19_En18
  input [18:0] Wgt_2_309, // sfix19_En18
  input [18:0] Wgt_2_310, // sfix19_En18
  input [18:0] Wgt_2_311, // sfix19_En18
  input [18:0] Wgt_2_312, // sfix19_En18
  input [18:0] Wgt_2_313, // sfix19_En18
  input [18:0] Wgt_2_314, // sfix19_En18
  input [18:0] Wgt_2_315, // sfix19_En18
  input [18:0] Wgt_2_316, // sfix19_En18
  input [18:0] Wgt_2_317, // sfix19_En18
  input [18:0] Wgt_2_318, // sfix19_En18
  input [18:0] Wgt_2_319, // sfix19_En18
  input [18:0] Wgt_2_320, // sfix19_En18
  input [18:0] Wgt_2_321, // sfix19_En18
  input [18:0] Wgt_2_322, // sfix19_En18
  input [18:0] Wgt_2_323, // sfix19_En18
  input [18:0] Wgt_2_324, // sfix19_En18
  input [18:0] Wgt_2_325, // sfix19_En18
  input [18:0] Wgt_2_326, // sfix19_En18
  input [18:0] Wgt_2_327, // sfix19_En18
  input [18:0] Wgt_2_328, // sfix19_En18
  input [18:0] Wgt_2_329, // sfix19_En18
  input [18:0] Wgt_2_330, // sfix19_En18
  input [18:0] Wgt_2_331, // sfix19_En18
  input [18:0] Wgt_2_332, // sfix19_En18
  input [18:0] Wgt_2_333, // sfix19_En18
  input [18:0] Wgt_2_334, // sfix19_En18
  input [18:0] Wgt_2_335, // sfix19_En18
  input [18:0] Wgt_2_336, // sfix19_En18
  input [18:0] Wgt_2_337, // sfix19_En18
  input [18:0] Wgt_2_338, // sfix19_En18
  input [18:0] Wgt_2_339, // sfix19_En18
  input [18:0] Wgt_2_340, // sfix19_En18
  input [18:0] Wgt_2_341, // sfix19_En18
  input [18:0] Wgt_2_342, // sfix19_En18
  input [18:0] Wgt_2_343, // sfix19_En18
  input [18:0] Wgt_2_344, // sfix19_En18
  input [18:0] Wgt_2_345, // sfix19_En18
  input [18:0] Wgt_2_346, // sfix19_En18
  input [18:0] Wgt_2_347, // sfix19_En18
  input [18:0] Wgt_2_348, // sfix19_En18
  input [18:0] Wgt_2_349, // sfix19_En18
  input [18:0] Wgt_2_350, // sfix19_En18
  input [18:0] Wgt_2_351, // sfix19_En18
  input [18:0] Wgt_2_352, // sfix19_En18
  input [18:0] Wgt_2_353, // sfix19_En18
  input [18:0] Wgt_2_354, // sfix19_En18
  input [18:0] Wgt_2_355, // sfix19_En18
  input [18:0] Wgt_2_356, // sfix19_En18
  input [18:0] Wgt_2_357, // sfix19_En18
  input [18:0] Wgt_2_358, // sfix19_En18
  input [18:0] Wgt_2_359, // sfix19_En18
  input [18:0] Wgt_2_360, // sfix19_En18
  input [18:0] Wgt_2_361, // sfix19_En18
  input [18:0] Wgt_2_362, // sfix19_En18
  input [18:0] Wgt_2_363, // sfix19_En18
  input [18:0] Wgt_2_364, // sfix19_En18
  input [18:0] Wgt_2_365, // sfix19_En18
  input [18:0] Wgt_2_366, // sfix19_En18
  input [18:0] Wgt_2_367, // sfix19_En18
  input [18:0] Wgt_2_368, // sfix19_En18
  input [18:0] Wgt_2_369, // sfix19_En18
  input [18:0] Wgt_2_370, // sfix19_En18
  input [18:0] Wgt_2_371, // sfix19_En18
  input [18:0] Wgt_2_372, // sfix19_En18
  input [18:0] Wgt_2_373, // sfix19_En18
  input [18:0] Wgt_2_374, // sfix19_En18
  input [18:0] Wgt_2_375, // sfix19_En18
  input [18:0] Wgt_2_376, // sfix19_En18
  input [18:0] Wgt_2_377, // sfix19_En18
  input [18:0] Wgt_2_378, // sfix19_En18
  input [18:0] Wgt_2_379, // sfix19_En18
  input [18:0] Wgt_2_380, // sfix19_En18
  input [18:0] Wgt_2_381, // sfix19_En18
  input [18:0] Wgt_2_382, // sfix19_En18
  input [18:0] Wgt_2_383, // sfix19_En18
  input [18:0] Wgt_2_384, // sfix19_En18
  input [18:0] Wgt_2_385, // sfix19_En18
  input [18:0] Wgt_2_386, // sfix19_En18
  input [18:0] Wgt_2_387, // sfix19_En18
  input [18:0] Wgt_2_388, // sfix19_En18
  input [18:0] Wgt_2_389, // sfix19_En18
  input [18:0] Wgt_2_390, // sfix19_En18
  input [18:0] Wgt_2_391, // sfix19_En18
  input [18:0] Wgt_2_392, // sfix19_En18
  input [18:0] Wgt_2_393, // sfix19_En18
  input [18:0] Wgt_2_394, // sfix19_En18
  input [18:0] Wgt_2_395, // sfix19_En18
  input [18:0] Wgt_2_396, // sfix19_En18
  input [18:0] Wgt_2_397, // sfix19_En18
  input [18:0] Wgt_2_398, // sfix19_En18
  input [18:0] Wgt_2_399, // sfix19_En18
  input [18:0] Wgt_2_400, // sfix19_En18
  input [18:0] Wgt_2_401, // sfix19_En18
  input [18:0] Wgt_2_402, // sfix19_En18
  input [18:0] Wgt_2_403, // sfix19_En18
  input [18:0] Wgt_2_404, // sfix19_En18
  input [18:0] Wgt_2_405, // sfix19_En18
  input [18:0] Wgt_2_406, // sfix19_En18
  input [18:0] Wgt_2_407, // sfix19_En18
  input [18:0] Wgt_2_408, // sfix19_En18
  input [18:0] Wgt_2_409, // sfix19_En18
  input [18:0] Wgt_2_410, // sfix19_En18
  input [18:0] Wgt_2_411, // sfix19_En18
  input [18:0] Wgt_2_412, // sfix19_En18
  input [18:0] Wgt_2_413, // sfix19_En18
  input [18:0] Wgt_2_414, // sfix19_En18
  input [18:0] Wgt_2_415, // sfix19_En18
  input [18:0] Wgt_2_416, // sfix19_En18
  input [18:0] Wgt_2_417, // sfix19_En18
  input [18:0] Wgt_2_418, // sfix19_En18
  input [18:0] Wgt_2_419, // sfix19_En18
  input [18:0] Wgt_2_420, // sfix19_En18
  input [18:0] Wgt_2_421, // sfix19_En18
  input [18:0] Wgt_2_422, // sfix19_En18
  input [18:0] Wgt_2_423, // sfix19_En18
  input [18:0] Wgt_2_424, // sfix19_En18
  input [18:0] Wgt_2_425, // sfix19_En18
  input [18:0] Wgt_2_426, // sfix19_En18
  input [18:0] Wgt_2_427, // sfix19_En18
  input [18:0] Wgt_2_428, // sfix19_En18
  input [18:0] Wgt_2_429, // sfix19_En18
  input [18:0] Wgt_2_430, // sfix19_En18
  input [18:0] Wgt_2_431, // sfix19_En18
  input [18:0] Wgt_2_432, // sfix19_En18
  input [18:0] Wgt_2_433, // sfix19_En18
  input [18:0] Wgt_2_434, // sfix19_En18
  input [18:0] Wgt_2_435, // sfix19_En18
  input [18:0] Wgt_2_436, // sfix19_En18
  input [18:0] Wgt_2_437, // sfix19_En18
  input [18:0] Wgt_2_438, // sfix19_En18
  input [18:0] Wgt_2_439, // sfix19_En18
  input [18:0] Wgt_2_440, // sfix19_En18
  input [18:0] Wgt_2_441, // sfix19_En18
  input [18:0] Wgt_2_442, // sfix19_En18
  input [18:0] Wgt_2_443, // sfix19_En18
  input [18:0] Wgt_2_444, // sfix19_En18
  input [18:0] Wgt_2_445, // sfix19_En18
  input [18:0] Wgt_2_446, // sfix19_En18
  input [18:0] Wgt_2_447, // sfix19_En18
  input [18:0] Wgt_2_448, // sfix19_En18
  input [18:0] Wgt_2_449, // sfix19_En18
  input [18:0] Wgt_2_450, // sfix19_En18
  input [18:0] Wgt_2_451, // sfix19_En18
  input [18:0] Wgt_2_452, // sfix19_En18
  input [18:0] Wgt_2_453, // sfix19_En18
  input [18:0] Wgt_2_454, // sfix19_En18
  input [18:0] Wgt_2_455, // sfix19_En18
  input [18:0] Wgt_2_456, // sfix19_En18
  input [18:0] Wgt_2_457, // sfix19_En18
  input [18:0] Wgt_2_458, // sfix19_En18
  input [18:0] Wgt_2_459, // sfix19_En18
  input [18:0] Wgt_2_460, // sfix19_En18
  input [18:0] Wgt_2_461, // sfix19_En18
  input [18:0] Wgt_2_462, // sfix19_En18
  input [18:0] Wgt_2_463, // sfix19_En18
  input [18:0] Wgt_2_464, // sfix19_En18
  input [18:0] Wgt_2_465, // sfix19_En18
  input [18:0] Wgt_2_466, // sfix19_En18
  input [18:0] Wgt_2_467, // sfix19_En18
  input [18:0] Wgt_2_468, // sfix19_En18
  input [18:0] Wgt_2_469, // sfix19_En18
  input [18:0] Wgt_2_470, // sfix19_En18
  input [18:0] Wgt_2_471, // sfix19_En18
  input [18:0] Wgt_2_472, // sfix19_En18
  input [18:0] Wgt_2_473, // sfix19_En18
  input [18:0] Wgt_2_474, // sfix19_En18
  input [18:0] Wgt_2_475, // sfix19_En18
  input [18:0] Wgt_2_476, // sfix19_En18
  input [18:0] Wgt_2_477, // sfix19_En18
  input [18:0] Wgt_2_478, // sfix19_En18
  input [18:0] Wgt_2_479, // sfix19_En18
  input [18:0] Wgt_2_480, // sfix19_En18
  input [18:0] Wgt_2_481, // sfix19_En18
  input [18:0] Wgt_2_482, // sfix19_En18
  input [18:0] Wgt_2_483, // sfix19_En18
  input [18:0] Wgt_2_484, // sfix19_En18
  input [18:0] Wgt_2_485, // sfix19_En18
  input [18:0] Wgt_2_486, // sfix19_En18
  input [18:0] Wgt_2_487, // sfix19_En18
  input [18:0] Wgt_2_488, // sfix19_En18
  input [18:0] Wgt_2_489, // sfix19_En18
  input [18:0] Wgt_2_490, // sfix19_En18
  input [18:0] Wgt_2_491, // sfix19_En18
  input [18:0] Wgt_2_492, // sfix19_En18
  input [18:0] Wgt_2_493, // sfix19_En18
  input [18:0] Wgt_2_494, // sfix19_En18
  input [18:0] Wgt_2_495, // sfix19_En18
  input [18:0] Wgt_2_496, // sfix19_En18
  input [18:0] Wgt_2_497, // sfix19_En18
  input [18:0] Wgt_2_498, // sfix19_En18
  input [18:0] Wgt_2_499, // sfix19_En18
  input [18:0] Wgt_2_500, // sfix19_En18
  input [18:0] Wgt_2_501, // sfix19_En18
  input [18:0] Wgt_2_502, // sfix19_En18
  input [18:0] Wgt_2_503, // sfix19_En18
  input [18:0] Wgt_2_504, // sfix19_En18
  input [18:0] Wgt_2_505, // sfix19_En18
  input [18:0] Wgt_2_506, // sfix19_En18
  input [18:0] Wgt_2_507, // sfix19_En18
  input [18:0] Wgt_2_508, // sfix19_En18
  input [18:0] Wgt_2_509, // sfix19_En18
  input [18:0] Wgt_2_510, // sfix19_En18
  input [18:0] Wgt_2_511, // sfix19_En18
  input [18:0] Wgt_2_512, // sfix19_En18
  input [18:0] Wgt_2_513, // sfix19_En18
  input [18:0] Wgt_2_514, // sfix19_En18
  input [18:0] Wgt_2_515, // sfix19_En18
  input [18:0] Wgt_2_516, // sfix19_En18
  input [18:0] Wgt_2_517, // sfix19_En18
  input [18:0] Wgt_2_518, // sfix19_En18
  input [18:0] Wgt_2_519, // sfix19_En18
  input [18:0] Wgt_2_520, // sfix19_En18
  input [18:0] Wgt_2_521, // sfix19_En18
  input [18:0] Wgt_2_522, // sfix19_En18
  input [18:0] Wgt_2_523, // sfix19_En18
  input [18:0] Wgt_2_524, // sfix19_En18
  input [18:0] Wgt_2_525, // sfix19_En18
  input [18:0] Wgt_2_526, // sfix19_En18
  input [18:0] Wgt_2_527, // sfix19_En18
  input [18:0] Wgt_2_528, // sfix19_En18
  input [18:0] Wgt_2_529, // sfix19_En18
  input [18:0] Wgt_2_530, // sfix19_En18
  input [18:0] Wgt_2_531, // sfix19_En18
  input [18:0] Wgt_2_532, // sfix19_En18
  input [18:0] Wgt_2_533, // sfix19_En18
  input [18:0] Wgt_2_534, // sfix19_En18
  input [18:0] Wgt_2_535, // sfix19_En18
  input [18:0] Wgt_2_536, // sfix19_En18
  input [18:0] Wgt_2_537, // sfix19_En18
  input [18:0] Wgt_2_538, // sfix19_En18
  input [18:0] Wgt_2_539, // sfix19_En18
  input [18:0] Wgt_2_540, // sfix19_En18
  input [18:0] Wgt_2_541, // sfix19_En18
  input [18:0] Wgt_2_542, // sfix19_En18
  input [18:0] Wgt_2_543, // sfix19_En18
  input [18:0] Wgt_2_544, // sfix19_En18
  input [18:0] Wgt_2_545, // sfix19_En18
  input [18:0] Wgt_2_546, // sfix19_En18
  input [18:0] Wgt_2_547, // sfix19_En18
  input [18:0] Wgt_2_548, // sfix19_En18
  input [18:0] Wgt_2_549, // sfix19_En18
  input [18:0] Wgt_2_550, // sfix19_En18
  input [18:0] Wgt_2_551, // sfix19_En18
  input [18:0] Wgt_2_552, // sfix19_En18
  input [18:0] Wgt_2_553, // sfix19_En18
  input [18:0] Wgt_2_554, // sfix19_En18
  input [18:0] Wgt_2_555, // sfix19_En18
  input [18:0] Wgt_2_556, // sfix19_En18
  input [18:0] Wgt_2_557, // sfix19_En18
  input [18:0] Wgt_2_558, // sfix19_En18
  input [18:0] Wgt_2_559, // sfix19_En18
  input [18:0] Wgt_2_560, // sfix19_En18
  input [18:0] Wgt_2_561, // sfix19_En18
  input [18:0] Wgt_2_562, // sfix19_En18
  input [18:0] Wgt_2_563, // sfix19_En18
  input [18:0] Wgt_2_564, // sfix19_En18
  input [18:0] Wgt_2_565, // sfix19_En18
  input [18:0] Wgt_2_566, // sfix19_En18
  input [18:0] Wgt_2_567, // sfix19_En18
  input [18:0] Wgt_2_568, // sfix19_En18
  input [18:0] Wgt_2_569, // sfix19_En18
  input [18:0] Wgt_2_570, // sfix19_En18
  input [18:0] Wgt_2_571, // sfix19_En18
  input [18:0] Wgt_2_572, // sfix19_En18
  input [18:0] Wgt_2_573, // sfix19_En18
  input [18:0] Wgt_2_574, // sfix19_En18
  input [18:0] Wgt_2_575, // sfix19_En18
  input [18:0] Wgt_2_576, // sfix19_En18
  input [18:0] Wgt_2_577, // sfix19_En18
  input [18:0] Wgt_2_578, // sfix19_En18
  input [18:0] Wgt_2_579, // sfix19_En18
  input [18:0] Wgt_2_580, // sfix19_En18
  input [18:0] Wgt_2_581, // sfix19_En18
  input [18:0] Wgt_2_582, // sfix19_En18
  input [18:0] Wgt_2_583, // sfix19_En18
  input [18:0] Wgt_2_584, // sfix19_En18
  input [18:0] Wgt_2_585, // sfix19_En18
  input [18:0] Wgt_2_586, // sfix19_En18
  input [18:0] Wgt_2_587, // sfix19_En18
  input [18:0] Wgt_2_588, // sfix19_En18
  input [18:0] Wgt_2_589, // sfix19_En18
  input [18:0] Wgt_2_590, // sfix19_En18
  input [18:0] Wgt_2_591, // sfix19_En18
  input [18:0] Wgt_2_592, // sfix19_En18
  input [18:0] Wgt_2_593, // sfix19_En18
  input [18:0] Wgt_2_594, // sfix19_En18
  input [18:0] Wgt_2_595, // sfix19_En18
  input [18:0] Wgt_2_596, // sfix19_En18
  input [18:0] Wgt_2_597, // sfix19_En18
  input [18:0] Wgt_2_598, // sfix19_En18
  input [18:0] Wgt_2_599, // sfix19_En18
  input [18:0] Wgt_2_600, // sfix19_En18
  input [18:0] Wgt_2_601, // sfix19_En18
  input [18:0] Wgt_2_602, // sfix19_En18
  input [18:0] Wgt_2_603, // sfix19_En18
  input [18:0] Wgt_2_604, // sfix19_En18
  input [18:0] Wgt_2_605, // sfix19_En18
  input [18:0] Wgt_2_606, // sfix19_En18
  input [18:0] Wgt_2_607, // sfix19_En18
  input [18:0] Wgt_2_608, // sfix19_En18
  input [18:0] Wgt_2_609, // sfix19_En18
  input [18:0] Wgt_2_610, // sfix19_En18
  input [18:0] Wgt_2_611, // sfix19_En18
  input [18:0] Wgt_2_612, // sfix19_En18
  input [18:0] Wgt_2_613, // sfix19_En18
  input [18:0] Wgt_2_614, // sfix19_En18
  input [18:0] Wgt_2_615, // sfix19_En18
  input [18:0] Wgt_2_616, // sfix19_En18
  input [18:0] Wgt_2_617, // sfix19_En18
  input [18:0] Wgt_2_618, // sfix19_En18
  input [18:0] Wgt_2_619, // sfix19_En18
  input [18:0] Wgt_2_620, // sfix19_En18
  input [18:0] Wgt_2_621, // sfix19_En18
  input [18:0] Wgt_2_622, // sfix19_En18
  input [18:0] Wgt_2_623, // sfix19_En18
  input [18:0] Wgt_2_624, // sfix19_En18
  input [18:0] Wgt_2_625, // sfix19_En18
  input [18:0] Wgt_2_626, // sfix19_En18
  input [18:0] Wgt_2_627, // sfix19_En18
  input [18:0] Wgt_2_628, // sfix19_En18
  input [18:0] Wgt_2_629, // sfix19_En18
  input [18:0] Wgt_2_630, // sfix19_En18
  input [18:0] Wgt_2_631, // sfix19_En18
  input [18:0] Wgt_2_632, // sfix19_En18
  input [18:0] Wgt_2_633, // sfix19_En18
  input [18:0] Wgt_2_634, // sfix19_En18
  input [18:0] Wgt_2_635, // sfix19_En18
  input [18:0] Wgt_2_636, // sfix19_En18
  input [18:0] Wgt_2_637, // sfix19_En18
  input [18:0] Wgt_2_638, // sfix19_En18
  input [18:0] Wgt_2_639, // sfix19_En18
  input [18:0] Wgt_2_640, // sfix19_En18
  input [18:0] Wgt_2_641, // sfix19_En18
  input [18:0] Wgt_2_642, // sfix19_En18
  input [18:0] Wgt_2_643, // sfix19_En18
  input [18:0] Wgt_2_644, // sfix19_En18
  input [18:0] Wgt_2_645, // sfix19_En18
  input [18:0] Wgt_2_646, // sfix19_En18
  input [18:0] Wgt_2_647, // sfix19_En18
  input [18:0] Wgt_2_648, // sfix19_En18
  input [18:0] Wgt_2_649, // sfix19_En18
  input [18:0] Wgt_2_650, // sfix19_En18
  input [18:0] Wgt_2_651, // sfix19_En18
  input [18:0] Wgt_2_652, // sfix19_En18
  input [18:0] Wgt_2_653, // sfix19_En18
  input [18:0] Wgt_2_654, // sfix19_En18
  input [18:0] Wgt_2_655, // sfix19_En18
  input [18:0] Wgt_2_656, // sfix19_En18
  input [18:0] Wgt_2_657, // sfix19_En18
  input [18:0] Wgt_2_658, // sfix19_En18
  input [18:0] Wgt_2_659, // sfix19_En18
  input [18:0] Wgt_2_660, // sfix19_En18
  input [18:0] Wgt_2_661, // sfix19_En18
  input [18:0] Wgt_2_662, // sfix19_En18
  input [18:0] Wgt_2_663, // sfix19_En18
  input [18:0] Wgt_2_664, // sfix19_En18
  input [18:0] Wgt_2_665, // sfix19_En18
  input [18:0] Wgt_2_666, // sfix19_En18
  input [18:0] Wgt_2_667, // sfix19_En18
  input [18:0] Wgt_2_668, // sfix19_En18
  input [18:0] Wgt_2_669, // sfix19_En18
  input [18:0] Wgt_2_670, // sfix19_En18
  input [18:0] Wgt_2_671, // sfix19_En18
  input [18:0] Wgt_2_672, // sfix19_En18
  input [18:0] Wgt_2_673, // sfix19_En18
  input [18:0] Wgt_2_674, // sfix19_En18
  input [18:0] Wgt_2_675, // sfix19_En18
  input [18:0] Wgt_2_676, // sfix19_En18
  input [18:0] Wgt_2_677, // sfix19_En18
  input [18:0] Wgt_2_678, // sfix19_En18
  input [18:0] Wgt_2_679, // sfix19_En18
  input [18:0] Wgt_2_680, // sfix19_En18
  input [18:0] Wgt_2_681, // sfix19_En18
  input [18:0] Wgt_2_682, // sfix19_En18
  input [18:0] Wgt_2_683, // sfix19_En18
  input [18:0] Wgt_2_684, // sfix19_En18
  input [18:0] Wgt_2_685, // sfix19_En18
  input [18:0] Wgt_2_686, // sfix19_En18
  input [18:0] Wgt_2_687, // sfix19_En18
  input [18:0] Wgt_2_688, // sfix19_En18
  input [18:0] Wgt_2_689, // sfix19_En18
  input [18:0] Wgt_2_690, // sfix19_En18
  input [18:0] Wgt_2_691, // sfix19_En18
  input [18:0] Wgt_2_692, // sfix19_En18
  input [18:0] Wgt_2_693, // sfix19_En18
  input [18:0] Wgt_2_694, // sfix19_En18
  input [18:0] Wgt_2_695, // sfix19_En18
  input [18:0] Wgt_2_696, // sfix19_En18
  input [18:0] Wgt_2_697, // sfix19_En18
  input [18:0] Wgt_2_698, // sfix19_En18
  input [18:0] Wgt_2_699, // sfix19_En18
  input [18:0] Wgt_2_700, // sfix19_En18
  input [18:0] Wgt_2_701, // sfix19_En18
  input [18:0] Wgt_2_702, // sfix19_En18
  input [18:0] Wgt_2_703, // sfix19_En18
  input [18:0] Wgt_2_704, // sfix19_En18
  input [18:0] Wgt_2_705, // sfix19_En18
  input [18:0] Wgt_2_706, // sfix19_En18
  input [18:0] Wgt_2_707, // sfix19_En18
  input [18:0] Wgt_2_708, // sfix19_En18
  input [18:0] Wgt_2_709, // sfix19_En18
  input [18:0] Wgt_2_710, // sfix19_En18
  input [18:0] Wgt_2_711, // sfix19_En18
  input [18:0] Wgt_2_712, // sfix19_En18
  input [18:0] Wgt_2_713, // sfix19_En18
  input [18:0] Wgt_2_714, // sfix19_En18
  input [18:0] Wgt_2_715, // sfix19_En18
  input [18:0] Wgt_2_716, // sfix19_En18
  input [18:0] Wgt_2_717, // sfix19_En18
  input [18:0] Wgt_2_718, // sfix19_En18
  input [18:0] Wgt_2_719, // sfix19_En18
  input [18:0] Wgt_2_720, // sfix19_En18
  input [18:0] Wgt_2_721, // sfix19_En18
  input [18:0] Wgt_2_722, // sfix19_En18
  input [18:0] Wgt_2_723, // sfix19_En18
  input [18:0] Wgt_2_724, // sfix19_En18
  input [18:0] Wgt_2_725, // sfix19_En18
  input [18:0] Wgt_2_726, // sfix19_En18
  input [18:0] Wgt_2_727, // sfix19_En18
  input [18:0] Wgt_2_728, // sfix19_En18
  input [18:0] Wgt_2_729, // sfix19_En18
  input [18:0] Wgt_2_730, // sfix19_En18
  input [18:0] Wgt_2_731, // sfix19_En18
  input [18:0] Wgt_2_732, // sfix19_En18
  input [18:0] Wgt_2_733, // sfix19_En18
  input [18:0] Wgt_2_734, // sfix19_En18
  input [18:0] Wgt_2_735, // sfix19_En18
  input [18:0] Wgt_2_736, // sfix19_En18
  input [18:0] Wgt_2_737, // sfix19_En18
  input [18:0] Wgt_2_738, // sfix19_En18
  input [18:0] Wgt_2_739, // sfix19_En18
  input [18:0] Wgt_2_740, // sfix19_En18
  input [18:0] Wgt_2_741, // sfix19_En18
  input [18:0] Wgt_2_742, // sfix19_En18
  input [18:0] Wgt_2_743, // sfix19_En18
  input [18:0] Wgt_2_744, // sfix19_En18
  input [18:0] Wgt_2_745, // sfix19_En18
  input [18:0] Wgt_2_746, // sfix19_En18
  input [18:0] Wgt_2_747, // sfix19_En18
  input [18:0] Wgt_2_748, // sfix19_En18
  input [18:0] Wgt_2_749, // sfix19_En18
  input [18:0] Wgt_2_750, // sfix19_En18
  input [18:0] Wgt_2_751, // sfix19_En18
  input [18:0] Wgt_2_752, // sfix19_En18
  input [18:0] Wgt_2_753, // sfix19_En18
  input [18:0] Wgt_2_754, // sfix19_En18
  input [18:0] Wgt_2_755, // sfix19_En18
  input [18:0] Wgt_2_756, // sfix19_En18
  input [18:0] Wgt_2_757, // sfix19_En18
  input [18:0] Wgt_2_758, // sfix19_En18
  input [18:0] Wgt_2_759, // sfix19_En18
  input [18:0] Wgt_2_760, // sfix19_En18
  input [18:0] Wgt_2_761, // sfix19_En18
  input [18:0] Wgt_2_762, // sfix19_En18
  input [18:0] Wgt_2_763, // sfix19_En18
  input [18:0] Wgt_2_764, // sfix19_En18
  input [18:0] Wgt_2_765, // sfix19_En18
  input [18:0] Wgt_2_766, // sfix19_En18
  input [18:0] Wgt_2_767, // sfix19_En18
  input [18:0] Wgt_2_768, // sfix19_En18
  input [18:0] Wgt_2_769, // sfix19_En18
  input [18:0] Wgt_2_770, // sfix19_En18
  input [18:0] Wgt_2_771, // sfix19_En18
  input [18:0] Wgt_2_772, // sfix19_En18
  input [18:0] Wgt_2_773, // sfix19_En18
  input [18:0] Wgt_2_774, // sfix19_En18
  input [18:0] Wgt_2_775, // sfix19_En18
  input [18:0] Wgt_2_776, // sfix19_En18
  input [18:0] Wgt_2_777, // sfix19_En18
  input [18:0] Wgt_2_778, // sfix19_En18
  input [18:0] Wgt_2_779, // sfix19_En18
  input [18:0] Wgt_2_780, // sfix19_En18
  input [18:0] Wgt_2_781, // sfix19_En18
  input [18:0] Wgt_2_782, // sfix19_En18
  input [18:0] Wgt_2_783, // sfix19_En18
  input [18:0] Wgt_2_784, // sfix19_En18
  input [18:0] Wgt_3_0, // sfix19_En18
  input [18:0] Wgt_3_1, // sfix19_En18
  input [18:0] Wgt_3_2, // sfix19_En18
  input [18:0] Wgt_3_3, // sfix19_En18
  input [18:0] Wgt_3_4, // sfix19_En18
  input [18:0] Wgt_3_5, // sfix19_En18
  input [18:0] Wgt_3_6, // sfix19_En18
  input [18:0] Wgt_3_7, // sfix19_En18
  input [18:0] Wgt_3_8, // sfix19_En18
  input [18:0] Wgt_3_9, // sfix19_En18
  input [18:0] Wgt_3_10, // sfix19_En18
  input [18:0] Wgt_3_11, // sfix19_En18
  input [18:0] Wgt_3_12, // sfix19_En18
  input [18:0] Wgt_3_13, // sfix19_En18
  input [18:0] Wgt_3_14, // sfix19_En18
  input [18:0] Wgt_3_15, // sfix19_En18
  input [18:0] Wgt_3_16, // sfix19_En18
  input [18:0] Wgt_3_17, // sfix19_En18
  input [18:0] Wgt_3_18, // sfix19_En18
  input [18:0] Wgt_3_19, // sfix19_En18
  input [18:0] Wgt_3_20, // sfix19_En18
  input [18:0] Wgt_3_21, // sfix19_En18
  input [18:0] Wgt_3_22, // sfix19_En18
  input [18:0] Wgt_3_23, // sfix19_En18
  input [18:0] Wgt_3_24, // sfix19_En18
  input [18:0] Wgt_3_25, // sfix19_En18
  input [18:0] Wgt_3_26, // sfix19_En18
  input [18:0] Wgt_3_27, // sfix19_En18
  input [18:0] Wgt_3_28, // sfix19_En18
  input [18:0] Wgt_3_29, // sfix19_En18
  input [18:0] Wgt_3_30, // sfix19_En18
  input [18:0] Wgt_3_31, // sfix19_En18
  input [18:0] Wgt_3_32, // sfix19_En18
  input [18:0] Wgt_3_33, // sfix19_En18
  input [18:0] Wgt_3_34, // sfix19_En18
  input [18:0] Wgt_3_35, // sfix19_En18
  input [18:0] Wgt_3_36, // sfix19_En18
  input [18:0] Wgt_3_37, // sfix19_En18
  input [18:0] Wgt_3_38, // sfix19_En18
  input [18:0] Wgt_3_39, // sfix19_En18
  input [18:0] Wgt_3_40, // sfix19_En18
  input [18:0] Wgt_3_41, // sfix19_En18
  input [18:0] Wgt_3_42, // sfix19_En18
  input [18:0] Wgt_3_43, // sfix19_En18
  input [18:0] Wgt_3_44, // sfix19_En18
  input [18:0] Wgt_3_45, // sfix19_En18
  input [18:0] Wgt_3_46, // sfix19_En18
  input [18:0] Wgt_3_47, // sfix19_En18
  input [18:0] Wgt_3_48, // sfix19_En18
  input [18:0] Wgt_3_49, // sfix19_En18
  input [18:0] Wgt_3_50, // sfix19_En18
  input [18:0] Wgt_3_51, // sfix19_En18
  input [18:0] Wgt_3_52, // sfix19_En18
  input [18:0] Wgt_3_53, // sfix19_En18
  input [18:0] Wgt_3_54, // sfix19_En18
  input [18:0] Wgt_3_55, // sfix19_En18
  input [18:0] Wgt_3_56, // sfix19_En18
  input [18:0] Wgt_3_57, // sfix19_En18
  input [18:0] Wgt_3_58, // sfix19_En18
  input [18:0] Wgt_3_59, // sfix19_En18
  input [18:0] Wgt_3_60, // sfix19_En18
  input [18:0] Wgt_3_61, // sfix19_En18
  input [18:0] Wgt_3_62, // sfix19_En18
  input [18:0] Wgt_3_63, // sfix19_En18
  input [18:0] Wgt_3_64, // sfix19_En18
  input [18:0] Wgt_3_65, // sfix19_En18
  input [18:0] Wgt_3_66, // sfix19_En18
  input [18:0] Wgt_3_67, // sfix19_En18
  input [18:0] Wgt_3_68, // sfix19_En18
  input [18:0] Wgt_3_69, // sfix19_En18
  input [18:0] Wgt_3_70, // sfix19_En18
  input [18:0] Wgt_3_71, // sfix19_En18
  input [18:0] Wgt_3_72, // sfix19_En18
  input [18:0] Wgt_3_73, // sfix19_En18
  input [18:0] Wgt_3_74, // sfix19_En18
  input [18:0] Wgt_3_75, // sfix19_En18
  input [18:0] Wgt_3_76, // sfix19_En18
  input [18:0] Wgt_3_77, // sfix19_En18
  input [18:0] Wgt_3_78, // sfix19_En18
  input [18:0] Wgt_3_79, // sfix19_En18
  input [18:0] Wgt_3_80, // sfix19_En18
  input [18:0] Wgt_3_81, // sfix19_En18
  input [18:0] Wgt_3_82, // sfix19_En18
  input [18:0] Wgt_3_83, // sfix19_En18
  input [18:0] Wgt_3_84, // sfix19_En18
  input [18:0] Wgt_3_85, // sfix19_En18
  input [18:0] Wgt_3_86, // sfix19_En18
  input [18:0] Wgt_3_87, // sfix19_En18
  input [18:0] Wgt_3_88, // sfix19_En18
  input [18:0] Wgt_3_89, // sfix19_En18
  input [18:0] Wgt_3_90, // sfix19_En18
  input [18:0] Wgt_3_91, // sfix19_En18
  input [18:0] Wgt_3_92, // sfix19_En18
  input [18:0] Wgt_3_93, // sfix19_En18
  input [18:0] Wgt_3_94, // sfix19_En18
  input [18:0] Wgt_3_95, // sfix19_En18
  input [18:0] Wgt_3_96, // sfix19_En18
  input [18:0] Wgt_3_97, // sfix19_En18
  input [18:0] Wgt_3_98, // sfix19_En18
  input [18:0] Wgt_3_99, // sfix19_En18
  input [18:0] Wgt_3_100, // sfix19_En18
  input [18:0] Wgt_3_101, // sfix19_En18
  input [18:0] Wgt_3_102, // sfix19_En18
  input [18:0] Wgt_3_103, // sfix19_En18
  input [18:0] Wgt_3_104, // sfix19_En18
  input [18:0] Wgt_3_105, // sfix19_En18
  input [18:0] Wgt_3_106, // sfix19_En18
  input [18:0] Wgt_3_107, // sfix19_En18
  input [18:0] Wgt_3_108, // sfix19_En18
  input [18:0] Wgt_3_109, // sfix19_En18
  input [18:0] Wgt_3_110, // sfix19_En18
  input [18:0] Wgt_3_111, // sfix19_En18
  input [18:0] Wgt_3_112, // sfix19_En18
  input [18:0] Wgt_3_113, // sfix19_En18
  input [18:0] Wgt_3_114, // sfix19_En18
  input [18:0] Wgt_3_115, // sfix19_En18
  input [18:0] Wgt_3_116, // sfix19_En18
  input [18:0] Wgt_3_117, // sfix19_En18
  input [18:0] Wgt_3_118, // sfix19_En18
  input [18:0] Wgt_3_119, // sfix19_En18
  input [18:0] Wgt_3_120, // sfix19_En18
  input [18:0] Wgt_3_121, // sfix19_En18
  input [18:0] Wgt_3_122, // sfix19_En18
  input [18:0] Wgt_3_123, // sfix19_En18
  input [18:0] Wgt_3_124, // sfix19_En18
  input [18:0] Wgt_3_125, // sfix19_En18
  input [18:0] Wgt_3_126, // sfix19_En18
  input [18:0] Wgt_3_127, // sfix19_En18
  input [18:0] Wgt_3_128, // sfix19_En18
  input [18:0] Wgt_3_129, // sfix19_En18
  input [18:0] Wgt_3_130, // sfix19_En18
  input [18:0] Wgt_3_131, // sfix19_En18
  input [18:0] Wgt_3_132, // sfix19_En18
  input [18:0] Wgt_3_133, // sfix19_En18
  input [18:0] Wgt_3_134, // sfix19_En18
  input [18:0] Wgt_3_135, // sfix19_En18
  input [18:0] Wgt_3_136, // sfix19_En18
  input [18:0] Wgt_3_137, // sfix19_En18
  input [18:0] Wgt_3_138, // sfix19_En18
  input [18:0] Wgt_3_139, // sfix19_En18
  input [18:0] Wgt_3_140, // sfix19_En18
  input [18:0] Wgt_3_141, // sfix19_En18
  input [18:0] Wgt_3_142, // sfix19_En18
  input [18:0] Wgt_3_143, // sfix19_En18
  input [18:0] Wgt_3_144, // sfix19_En18
  input [18:0] Wgt_3_145, // sfix19_En18
  input [18:0] Wgt_3_146, // sfix19_En18
  input [18:0] Wgt_3_147, // sfix19_En18
  input [18:0] Wgt_3_148, // sfix19_En18
  input [18:0] Wgt_3_149, // sfix19_En18
  input [18:0] Wgt_3_150, // sfix19_En18
  input [18:0] Wgt_3_151, // sfix19_En18
  input [18:0] Wgt_3_152, // sfix19_En18
  input [18:0] Wgt_3_153, // sfix19_En18
  input [18:0] Wgt_3_154, // sfix19_En18
  input [18:0] Wgt_3_155, // sfix19_En18
  input [18:0] Wgt_3_156, // sfix19_En18
  input [18:0] Wgt_3_157, // sfix19_En18
  input [18:0] Wgt_3_158, // sfix19_En18
  input [18:0] Wgt_3_159, // sfix19_En18
  input [18:0] Wgt_3_160, // sfix19_En18
  input [18:0] Wgt_3_161, // sfix19_En18
  input [18:0] Wgt_3_162, // sfix19_En18
  input [18:0] Wgt_3_163, // sfix19_En18
  input [18:0] Wgt_3_164, // sfix19_En18
  input [18:0] Wgt_3_165, // sfix19_En18
  input [18:0] Wgt_3_166, // sfix19_En18
  input [18:0] Wgt_3_167, // sfix19_En18
  input [18:0] Wgt_3_168, // sfix19_En18
  input [18:0] Wgt_3_169, // sfix19_En18
  input [18:0] Wgt_3_170, // sfix19_En18
  input [18:0] Wgt_3_171, // sfix19_En18
  input [18:0] Wgt_3_172, // sfix19_En18
  input [18:0] Wgt_3_173, // sfix19_En18
  input [18:0] Wgt_3_174, // sfix19_En18
  input [18:0] Wgt_3_175, // sfix19_En18
  input [18:0] Wgt_3_176, // sfix19_En18
  input [18:0] Wgt_3_177, // sfix19_En18
  input [18:0] Wgt_3_178, // sfix19_En18
  input [18:0] Wgt_3_179, // sfix19_En18
  input [18:0] Wgt_3_180, // sfix19_En18
  input [18:0] Wgt_3_181, // sfix19_En18
  input [18:0] Wgt_3_182, // sfix19_En18
  input [18:0] Wgt_3_183, // sfix19_En18
  input [18:0] Wgt_3_184, // sfix19_En18
  input [18:0] Wgt_3_185, // sfix19_En18
  input [18:0] Wgt_3_186, // sfix19_En18
  input [18:0] Wgt_3_187, // sfix19_En18
  input [18:0] Wgt_3_188, // sfix19_En18
  input [18:0] Wgt_3_189, // sfix19_En18
  input [18:0] Wgt_3_190, // sfix19_En18
  input [18:0] Wgt_3_191, // sfix19_En18
  input [18:0] Wgt_3_192, // sfix19_En18
  input [18:0] Wgt_3_193, // sfix19_En18
  input [18:0] Wgt_3_194, // sfix19_En18
  input [18:0] Wgt_3_195, // sfix19_En18
  input [18:0] Wgt_3_196, // sfix19_En18
  input [18:0] Wgt_3_197, // sfix19_En18
  input [18:0] Wgt_3_198, // sfix19_En18
  input [18:0] Wgt_3_199, // sfix19_En18
  input [18:0] Wgt_3_200, // sfix19_En18
  input [18:0] Wgt_3_201, // sfix19_En18
  input [18:0] Wgt_3_202, // sfix19_En18
  input [18:0] Wgt_3_203, // sfix19_En18
  input [18:0] Wgt_3_204, // sfix19_En18
  input [18:0] Wgt_3_205, // sfix19_En18
  input [18:0] Wgt_3_206, // sfix19_En18
  input [18:0] Wgt_3_207, // sfix19_En18
  input [18:0] Wgt_3_208, // sfix19_En18
  input [18:0] Wgt_3_209, // sfix19_En18
  input [18:0] Wgt_3_210, // sfix19_En18
  input [18:0] Wgt_3_211, // sfix19_En18
  input [18:0] Wgt_3_212, // sfix19_En18
  input [18:0] Wgt_3_213, // sfix19_En18
  input [18:0] Wgt_3_214, // sfix19_En18
  input [18:0] Wgt_3_215, // sfix19_En18
  input [18:0] Wgt_3_216, // sfix19_En18
  input [18:0] Wgt_3_217, // sfix19_En18
  input [18:0] Wgt_3_218, // sfix19_En18
  input [18:0] Wgt_3_219, // sfix19_En18
  input [18:0] Wgt_3_220, // sfix19_En18
  input [18:0] Wgt_3_221, // sfix19_En18
  input [18:0] Wgt_3_222, // sfix19_En18
  input [18:0] Wgt_3_223, // sfix19_En18
  input [18:0] Wgt_3_224, // sfix19_En18
  input [18:0] Wgt_3_225, // sfix19_En18
  input [18:0] Wgt_3_226, // sfix19_En18
  input [18:0] Wgt_3_227, // sfix19_En18
  input [18:0] Wgt_3_228, // sfix19_En18
  input [18:0] Wgt_3_229, // sfix19_En18
  input [18:0] Wgt_3_230, // sfix19_En18
  input [18:0] Wgt_3_231, // sfix19_En18
  input [18:0] Wgt_3_232, // sfix19_En18
  input [18:0] Wgt_3_233, // sfix19_En18
  input [18:0] Wgt_3_234, // sfix19_En18
  input [18:0] Wgt_3_235, // sfix19_En18
  input [18:0] Wgt_3_236, // sfix19_En18
  input [18:0] Wgt_3_237, // sfix19_En18
  input [18:0] Wgt_3_238, // sfix19_En18
  input [18:0] Wgt_3_239, // sfix19_En18
  input [18:0] Wgt_3_240, // sfix19_En18
  input [18:0] Wgt_3_241, // sfix19_En18
  input [18:0] Wgt_3_242, // sfix19_En18
  input [18:0] Wgt_3_243, // sfix19_En18
  input [18:0] Wgt_3_244, // sfix19_En18
  input [18:0] Wgt_3_245, // sfix19_En18
  input [18:0] Wgt_3_246, // sfix19_En18
  input [18:0] Wgt_3_247, // sfix19_En18
  input [18:0] Wgt_3_248, // sfix19_En18
  input [18:0] Wgt_3_249, // sfix19_En18
  input [18:0] Wgt_3_250, // sfix19_En18
  input [18:0] Wgt_3_251, // sfix19_En18
  input [18:0] Wgt_3_252, // sfix19_En18
  input [18:0] Wgt_3_253, // sfix19_En18
  input [18:0] Wgt_3_254, // sfix19_En18
  input [18:0] Wgt_3_255, // sfix19_En18
  input [18:0] Wgt_3_256, // sfix19_En18
  input [18:0] Wgt_3_257, // sfix19_En18
  input [18:0] Wgt_3_258, // sfix19_En18
  input [18:0] Wgt_3_259, // sfix19_En18
  input [18:0] Wgt_3_260, // sfix19_En18
  input [18:0] Wgt_3_261, // sfix19_En18
  input [18:0] Wgt_3_262, // sfix19_En18
  input [18:0] Wgt_3_263, // sfix19_En18
  input [18:0] Wgt_3_264, // sfix19_En18
  input [18:0] Wgt_3_265, // sfix19_En18
  input [18:0] Wgt_3_266, // sfix19_En18
  input [18:0] Wgt_3_267, // sfix19_En18
  input [18:0] Wgt_3_268, // sfix19_En18
  input [18:0] Wgt_3_269, // sfix19_En18
  input [18:0] Wgt_3_270, // sfix19_En18
  input [18:0] Wgt_3_271, // sfix19_En18
  input [18:0] Wgt_3_272, // sfix19_En18
  input [18:0] Wgt_3_273, // sfix19_En18
  input [18:0] Wgt_3_274, // sfix19_En18
  input [18:0] Wgt_3_275, // sfix19_En18
  input [18:0] Wgt_3_276, // sfix19_En18
  input [18:0] Wgt_3_277, // sfix19_En18
  input [18:0] Wgt_3_278, // sfix19_En18
  input [18:0] Wgt_3_279, // sfix19_En18
  input [18:0] Wgt_3_280, // sfix19_En18
  input [18:0] Wgt_3_281, // sfix19_En18
  input [18:0] Wgt_3_282, // sfix19_En18
  input [18:0] Wgt_3_283, // sfix19_En18
  input [18:0] Wgt_3_284, // sfix19_En18
  input [18:0] Wgt_3_285, // sfix19_En18
  input [18:0] Wgt_3_286, // sfix19_En18
  input [18:0] Wgt_3_287, // sfix19_En18
  input [18:0] Wgt_3_288, // sfix19_En18
  input [18:0] Wgt_3_289, // sfix19_En18
  input [18:0] Wgt_3_290, // sfix19_En18
  input [18:0] Wgt_3_291, // sfix19_En18
  input [18:0] Wgt_3_292, // sfix19_En18
  input [18:0] Wgt_3_293, // sfix19_En18
  input [18:0] Wgt_3_294, // sfix19_En18
  input [18:0] Wgt_3_295, // sfix19_En18
  input [18:0] Wgt_3_296, // sfix19_En18
  input [18:0] Wgt_3_297, // sfix19_En18
  input [18:0] Wgt_3_298, // sfix19_En18
  input [18:0] Wgt_3_299, // sfix19_En18
  input [18:0] Wgt_3_300, // sfix19_En18
  input [18:0] Wgt_3_301, // sfix19_En18
  input [18:0] Wgt_3_302, // sfix19_En18
  input [18:0] Wgt_3_303, // sfix19_En18
  input [18:0] Wgt_3_304, // sfix19_En18
  input [18:0] Wgt_3_305, // sfix19_En18
  input [18:0] Wgt_3_306, // sfix19_En18
  input [18:0] Wgt_3_307, // sfix19_En18
  input [18:0] Wgt_3_308, // sfix19_En18
  input [18:0] Wgt_3_309, // sfix19_En18
  input [18:0] Wgt_3_310, // sfix19_En18
  input [18:0] Wgt_3_311, // sfix19_En18
  input [18:0] Wgt_3_312, // sfix19_En18
  input [18:0] Wgt_3_313, // sfix19_En18
  input [18:0] Wgt_3_314, // sfix19_En18
  input [18:0] Wgt_3_315, // sfix19_En18
  input [18:0] Wgt_3_316, // sfix19_En18
  input [18:0] Wgt_3_317, // sfix19_En18
  input [18:0] Wgt_3_318, // sfix19_En18
  input [18:0] Wgt_3_319, // sfix19_En18
  input [18:0] Wgt_3_320, // sfix19_En18
  input [18:0] Wgt_3_321, // sfix19_En18
  input [18:0] Wgt_3_322, // sfix19_En18
  input [18:0] Wgt_3_323, // sfix19_En18
  input [18:0] Wgt_3_324, // sfix19_En18
  input [18:0] Wgt_3_325, // sfix19_En18
  input [18:0] Wgt_3_326, // sfix19_En18
  input [18:0] Wgt_3_327, // sfix19_En18
  input [18:0] Wgt_3_328, // sfix19_En18
  input [18:0] Wgt_3_329, // sfix19_En18
  input [18:0] Wgt_3_330, // sfix19_En18
  input [18:0] Wgt_3_331, // sfix19_En18
  input [18:0] Wgt_3_332, // sfix19_En18
  input [18:0] Wgt_3_333, // sfix19_En18
  input [18:0] Wgt_3_334, // sfix19_En18
  input [18:0] Wgt_3_335, // sfix19_En18
  input [18:0] Wgt_3_336, // sfix19_En18
  input [18:0] Wgt_3_337, // sfix19_En18
  input [18:0] Wgt_3_338, // sfix19_En18
  input [18:0] Wgt_3_339, // sfix19_En18
  input [18:0] Wgt_3_340, // sfix19_En18
  input [18:0] Wgt_3_341, // sfix19_En18
  input [18:0] Wgt_3_342, // sfix19_En18
  input [18:0] Wgt_3_343, // sfix19_En18
  input [18:0] Wgt_3_344, // sfix19_En18
  input [18:0] Wgt_3_345, // sfix19_En18
  input [18:0] Wgt_3_346, // sfix19_En18
  input [18:0] Wgt_3_347, // sfix19_En18
  input [18:0] Wgt_3_348, // sfix19_En18
  input [18:0] Wgt_3_349, // sfix19_En18
  input [18:0] Wgt_3_350, // sfix19_En18
  input [18:0] Wgt_3_351, // sfix19_En18
  input [18:0] Wgt_3_352, // sfix19_En18
  input [18:0] Wgt_3_353, // sfix19_En18
  input [18:0] Wgt_3_354, // sfix19_En18
  input [18:0] Wgt_3_355, // sfix19_En18
  input [18:0] Wgt_3_356, // sfix19_En18
  input [18:0] Wgt_3_357, // sfix19_En18
  input [18:0] Wgt_3_358, // sfix19_En18
  input [18:0] Wgt_3_359, // sfix19_En18
  input [18:0] Wgt_3_360, // sfix19_En18
  input [18:0] Wgt_3_361, // sfix19_En18
  input [18:0] Wgt_3_362, // sfix19_En18
  input [18:0] Wgt_3_363, // sfix19_En18
  input [18:0] Wgt_3_364, // sfix19_En18
  input [18:0] Wgt_3_365, // sfix19_En18
  input [18:0] Wgt_3_366, // sfix19_En18
  input [18:0] Wgt_3_367, // sfix19_En18
  input [18:0] Wgt_3_368, // sfix19_En18
  input [18:0] Wgt_3_369, // sfix19_En18
  input [18:0] Wgt_3_370, // sfix19_En18
  input [18:0] Wgt_3_371, // sfix19_En18
  input [18:0] Wgt_3_372, // sfix19_En18
  input [18:0] Wgt_3_373, // sfix19_En18
  input [18:0] Wgt_3_374, // sfix19_En18
  input [18:0] Wgt_3_375, // sfix19_En18
  input [18:0] Wgt_3_376, // sfix19_En18
  input [18:0] Wgt_3_377, // sfix19_En18
  input [18:0] Wgt_3_378, // sfix19_En18
  input [18:0] Wgt_3_379, // sfix19_En18
  input [18:0] Wgt_3_380, // sfix19_En18
  input [18:0] Wgt_3_381, // sfix19_En18
  input [18:0] Wgt_3_382, // sfix19_En18
  input [18:0] Wgt_3_383, // sfix19_En18
  input [18:0] Wgt_3_384, // sfix19_En18
  input [18:0] Wgt_3_385, // sfix19_En18
  input [18:0] Wgt_3_386, // sfix19_En18
  input [18:0] Wgt_3_387, // sfix19_En18
  input [18:0] Wgt_3_388, // sfix19_En18
  input [18:0] Wgt_3_389, // sfix19_En18
  input [18:0] Wgt_3_390, // sfix19_En18
  input [18:0] Wgt_3_391, // sfix19_En18
  input [18:0] Wgt_3_392, // sfix19_En18
  input [18:0] Wgt_3_393, // sfix19_En18
  input [18:0] Wgt_3_394, // sfix19_En18
  input [18:0] Wgt_3_395, // sfix19_En18
  input [18:0] Wgt_3_396, // sfix19_En18
  input [18:0] Wgt_3_397, // sfix19_En18
  input [18:0] Wgt_3_398, // sfix19_En18
  input [18:0] Wgt_3_399, // sfix19_En18
  input [18:0] Wgt_3_400, // sfix19_En18
  input [18:0] Wgt_3_401, // sfix19_En18
  input [18:0] Wgt_3_402, // sfix19_En18
  input [18:0] Wgt_3_403, // sfix19_En18
  input [18:0] Wgt_3_404, // sfix19_En18
  input [18:0] Wgt_3_405, // sfix19_En18
  input [18:0] Wgt_3_406, // sfix19_En18
  input [18:0] Wgt_3_407, // sfix19_En18
  input [18:0] Wgt_3_408, // sfix19_En18
  input [18:0] Wgt_3_409, // sfix19_En18
  input [18:0] Wgt_3_410, // sfix19_En18
  input [18:0] Wgt_3_411, // sfix19_En18
  input [18:0] Wgt_3_412, // sfix19_En18
  input [18:0] Wgt_3_413, // sfix19_En18
  input [18:0] Wgt_3_414, // sfix19_En18
  input [18:0] Wgt_3_415, // sfix19_En18
  input [18:0] Wgt_3_416, // sfix19_En18
  input [18:0] Wgt_3_417, // sfix19_En18
  input [18:0] Wgt_3_418, // sfix19_En18
  input [18:0] Wgt_3_419, // sfix19_En18
  input [18:0] Wgt_3_420, // sfix19_En18
  input [18:0] Wgt_3_421, // sfix19_En18
  input [18:0] Wgt_3_422, // sfix19_En18
  input [18:0] Wgt_3_423, // sfix19_En18
  input [18:0] Wgt_3_424, // sfix19_En18
  input [18:0] Wgt_3_425, // sfix19_En18
  input [18:0] Wgt_3_426, // sfix19_En18
  input [18:0] Wgt_3_427, // sfix19_En18
  input [18:0] Wgt_3_428, // sfix19_En18
  input [18:0] Wgt_3_429, // sfix19_En18
  input [18:0] Wgt_3_430, // sfix19_En18
  input [18:0] Wgt_3_431, // sfix19_En18
  input [18:0] Wgt_3_432, // sfix19_En18
  input [18:0] Wgt_3_433, // sfix19_En18
  input [18:0] Wgt_3_434, // sfix19_En18
  input [18:0] Wgt_3_435, // sfix19_En18
  input [18:0] Wgt_3_436, // sfix19_En18
  input [18:0] Wgt_3_437, // sfix19_En18
  input [18:0] Wgt_3_438, // sfix19_En18
  input [18:0] Wgt_3_439, // sfix19_En18
  input [18:0] Wgt_3_440, // sfix19_En18
  input [18:0] Wgt_3_441, // sfix19_En18
  input [18:0] Wgt_3_442, // sfix19_En18
  input [18:0] Wgt_3_443, // sfix19_En18
  input [18:0] Wgt_3_444, // sfix19_En18
  input [18:0] Wgt_3_445, // sfix19_En18
  input [18:0] Wgt_3_446, // sfix19_En18
  input [18:0] Wgt_3_447, // sfix19_En18
  input [18:0] Wgt_3_448, // sfix19_En18
  input [18:0] Wgt_3_449, // sfix19_En18
  input [18:0] Wgt_3_450, // sfix19_En18
  input [18:0] Wgt_3_451, // sfix19_En18
  input [18:0] Wgt_3_452, // sfix19_En18
  input [18:0] Wgt_3_453, // sfix19_En18
  input [18:0] Wgt_3_454, // sfix19_En18
  input [18:0] Wgt_3_455, // sfix19_En18
  input [18:0] Wgt_3_456, // sfix19_En18
  input [18:0] Wgt_3_457, // sfix19_En18
  input [18:0] Wgt_3_458, // sfix19_En18
  input [18:0] Wgt_3_459, // sfix19_En18
  input [18:0] Wgt_3_460, // sfix19_En18
  input [18:0] Wgt_3_461, // sfix19_En18
  input [18:0] Wgt_3_462, // sfix19_En18
  input [18:0] Wgt_3_463, // sfix19_En18
  input [18:0] Wgt_3_464, // sfix19_En18
  input [18:0] Wgt_3_465, // sfix19_En18
  input [18:0] Wgt_3_466, // sfix19_En18
  input [18:0] Wgt_3_467, // sfix19_En18
  input [18:0] Wgt_3_468, // sfix19_En18
  input [18:0] Wgt_3_469, // sfix19_En18
  input [18:0] Wgt_3_470, // sfix19_En18
  input [18:0] Wgt_3_471, // sfix19_En18
  input [18:0] Wgt_3_472, // sfix19_En18
  input [18:0] Wgt_3_473, // sfix19_En18
  input [18:0] Wgt_3_474, // sfix19_En18
  input [18:0] Wgt_3_475, // sfix19_En18
  input [18:0] Wgt_3_476, // sfix19_En18
  input [18:0] Wgt_3_477, // sfix19_En18
  input [18:0] Wgt_3_478, // sfix19_En18
  input [18:0] Wgt_3_479, // sfix19_En18
  input [18:0] Wgt_3_480, // sfix19_En18
  input [18:0] Wgt_3_481, // sfix19_En18
  input [18:0] Wgt_3_482, // sfix19_En18
  input [18:0] Wgt_3_483, // sfix19_En18
  input [18:0] Wgt_3_484, // sfix19_En18
  input [18:0] Wgt_3_485, // sfix19_En18
  input [18:0] Wgt_3_486, // sfix19_En18
  input [18:0] Wgt_3_487, // sfix19_En18
  input [18:0] Wgt_3_488, // sfix19_En18
  input [18:0] Wgt_3_489, // sfix19_En18
  input [18:0] Wgt_3_490, // sfix19_En18
  input [18:0] Wgt_3_491, // sfix19_En18
  input [18:0] Wgt_3_492, // sfix19_En18
  input [18:0] Wgt_3_493, // sfix19_En18
  input [18:0] Wgt_3_494, // sfix19_En18
  input [18:0] Wgt_3_495, // sfix19_En18
  input [18:0] Wgt_3_496, // sfix19_En18
  input [18:0] Wgt_3_497, // sfix19_En18
  input [18:0] Wgt_3_498, // sfix19_En18
  input [18:0] Wgt_3_499, // sfix19_En18
  input [18:0] Wgt_3_500, // sfix19_En18
  input [18:0] Wgt_3_501, // sfix19_En18
  input [18:0] Wgt_3_502, // sfix19_En18
  input [18:0] Wgt_3_503, // sfix19_En18
  input [18:0] Wgt_3_504, // sfix19_En18
  input [18:0] Wgt_3_505, // sfix19_En18
  input [18:0] Wgt_3_506, // sfix19_En18
  input [18:0] Wgt_3_507, // sfix19_En18
  input [18:0] Wgt_3_508, // sfix19_En18
  input [18:0] Wgt_3_509, // sfix19_En18
  input [18:0] Wgt_3_510, // sfix19_En18
  input [18:0] Wgt_3_511, // sfix19_En18
  input [18:0] Wgt_3_512, // sfix19_En18
  input [18:0] Wgt_3_513, // sfix19_En18
  input [18:0] Wgt_3_514, // sfix19_En18
  input [18:0] Wgt_3_515, // sfix19_En18
  input [18:0] Wgt_3_516, // sfix19_En18
  input [18:0] Wgt_3_517, // sfix19_En18
  input [18:0] Wgt_3_518, // sfix19_En18
  input [18:0] Wgt_3_519, // sfix19_En18
  input [18:0] Wgt_3_520, // sfix19_En18
  input [18:0] Wgt_3_521, // sfix19_En18
  input [18:0] Wgt_3_522, // sfix19_En18
  input [18:0] Wgt_3_523, // sfix19_En18
  input [18:0] Wgt_3_524, // sfix19_En18
  input [18:0] Wgt_3_525, // sfix19_En18
  input [18:0] Wgt_3_526, // sfix19_En18
  input [18:0] Wgt_3_527, // sfix19_En18
  input [18:0] Wgt_3_528, // sfix19_En18
  input [18:0] Wgt_3_529, // sfix19_En18
  input [18:0] Wgt_3_530, // sfix19_En18
  input [18:0] Wgt_3_531, // sfix19_En18
  input [18:0] Wgt_3_532, // sfix19_En18
  input [18:0] Wgt_3_533, // sfix19_En18
  input [18:0] Wgt_3_534, // sfix19_En18
  input [18:0] Wgt_3_535, // sfix19_En18
  input [18:0] Wgt_3_536, // sfix19_En18
  input [18:0] Wgt_3_537, // sfix19_En18
  input [18:0] Wgt_3_538, // sfix19_En18
  input [18:0] Wgt_3_539, // sfix19_En18
  input [18:0] Wgt_3_540, // sfix19_En18
  input [18:0] Wgt_3_541, // sfix19_En18
  input [18:0] Wgt_3_542, // sfix19_En18
  input [18:0] Wgt_3_543, // sfix19_En18
  input [18:0] Wgt_3_544, // sfix19_En18
  input [18:0] Wgt_3_545, // sfix19_En18
  input [18:0] Wgt_3_546, // sfix19_En18
  input [18:0] Wgt_3_547, // sfix19_En18
  input [18:0] Wgt_3_548, // sfix19_En18
  input [18:0] Wgt_3_549, // sfix19_En18
  input [18:0] Wgt_3_550, // sfix19_En18
  input [18:0] Wgt_3_551, // sfix19_En18
  input [18:0] Wgt_3_552, // sfix19_En18
  input [18:0] Wgt_3_553, // sfix19_En18
  input [18:0] Wgt_3_554, // sfix19_En18
  input [18:0] Wgt_3_555, // sfix19_En18
  input [18:0] Wgt_3_556, // sfix19_En18
  input [18:0] Wgt_3_557, // sfix19_En18
  input [18:0] Wgt_3_558, // sfix19_En18
  input [18:0] Wgt_3_559, // sfix19_En18
  input [18:0] Wgt_3_560, // sfix19_En18
  input [18:0] Wgt_3_561, // sfix19_En18
  input [18:0] Wgt_3_562, // sfix19_En18
  input [18:0] Wgt_3_563, // sfix19_En18
  input [18:0] Wgt_3_564, // sfix19_En18
  input [18:0] Wgt_3_565, // sfix19_En18
  input [18:0] Wgt_3_566, // sfix19_En18
  input [18:0] Wgt_3_567, // sfix19_En18
  input [18:0] Wgt_3_568, // sfix19_En18
  input [18:0] Wgt_3_569, // sfix19_En18
  input [18:0] Wgt_3_570, // sfix19_En18
  input [18:0] Wgt_3_571, // sfix19_En18
  input [18:0] Wgt_3_572, // sfix19_En18
  input [18:0] Wgt_3_573, // sfix19_En18
  input [18:0] Wgt_3_574, // sfix19_En18
  input [18:0] Wgt_3_575, // sfix19_En18
  input [18:0] Wgt_3_576, // sfix19_En18
  input [18:0] Wgt_3_577, // sfix19_En18
  input [18:0] Wgt_3_578, // sfix19_En18
  input [18:0] Wgt_3_579, // sfix19_En18
  input [18:0] Wgt_3_580, // sfix19_En18
  input [18:0] Wgt_3_581, // sfix19_En18
  input [18:0] Wgt_3_582, // sfix19_En18
  input [18:0] Wgt_3_583, // sfix19_En18
  input [18:0] Wgt_3_584, // sfix19_En18
  input [18:0] Wgt_3_585, // sfix19_En18
  input [18:0] Wgt_3_586, // sfix19_En18
  input [18:0] Wgt_3_587, // sfix19_En18
  input [18:0] Wgt_3_588, // sfix19_En18
  input [18:0] Wgt_3_589, // sfix19_En18
  input [18:0] Wgt_3_590, // sfix19_En18
  input [18:0] Wgt_3_591, // sfix19_En18
  input [18:0] Wgt_3_592, // sfix19_En18
  input [18:0] Wgt_3_593, // sfix19_En18
  input [18:0] Wgt_3_594, // sfix19_En18
  input [18:0] Wgt_3_595, // sfix19_En18
  input [18:0] Wgt_3_596, // sfix19_En18
  input [18:0] Wgt_3_597, // sfix19_En18
  input [18:0] Wgt_3_598, // sfix19_En18
  input [18:0] Wgt_3_599, // sfix19_En18
  input [18:0] Wgt_3_600, // sfix19_En18
  input [18:0] Wgt_3_601, // sfix19_En18
  input [18:0] Wgt_3_602, // sfix19_En18
  input [18:0] Wgt_3_603, // sfix19_En18
  input [18:0] Wgt_3_604, // sfix19_En18
  input [18:0] Wgt_3_605, // sfix19_En18
  input [18:0] Wgt_3_606, // sfix19_En18
  input [18:0] Wgt_3_607, // sfix19_En18
  input [18:0] Wgt_3_608, // sfix19_En18
  input [18:0] Wgt_3_609, // sfix19_En18
  input [18:0] Wgt_3_610, // sfix19_En18
  input [18:0] Wgt_3_611, // sfix19_En18
  input [18:0] Wgt_3_612, // sfix19_En18
  input [18:0] Wgt_3_613, // sfix19_En18
  input [18:0] Wgt_3_614, // sfix19_En18
  input [18:0] Wgt_3_615, // sfix19_En18
  input [18:0] Wgt_3_616, // sfix19_En18
  input [18:0] Wgt_3_617, // sfix19_En18
  input [18:0] Wgt_3_618, // sfix19_En18
  input [18:0] Wgt_3_619, // sfix19_En18
  input [18:0] Wgt_3_620, // sfix19_En18
  input [18:0] Wgt_3_621, // sfix19_En18
  input [18:0] Wgt_3_622, // sfix19_En18
  input [18:0] Wgt_3_623, // sfix19_En18
  input [18:0] Wgt_3_624, // sfix19_En18
  input [18:0] Wgt_3_625, // sfix19_En18
  input [18:0] Wgt_3_626, // sfix19_En18
  input [18:0] Wgt_3_627, // sfix19_En18
  input [18:0] Wgt_3_628, // sfix19_En18
  input [18:0] Wgt_3_629, // sfix19_En18
  input [18:0] Wgt_3_630, // sfix19_En18
  input [18:0] Wgt_3_631, // sfix19_En18
  input [18:0] Wgt_3_632, // sfix19_En18
  input [18:0] Wgt_3_633, // sfix19_En18
  input [18:0] Wgt_3_634, // sfix19_En18
  input [18:0] Wgt_3_635, // sfix19_En18
  input [18:0] Wgt_3_636, // sfix19_En18
  input [18:0] Wgt_3_637, // sfix19_En18
  input [18:0] Wgt_3_638, // sfix19_En18
  input [18:0] Wgt_3_639, // sfix19_En18
  input [18:0] Wgt_3_640, // sfix19_En18
  input [18:0] Wgt_3_641, // sfix19_En18
  input [18:0] Wgt_3_642, // sfix19_En18
  input [18:0] Wgt_3_643, // sfix19_En18
  input [18:0] Wgt_3_644, // sfix19_En18
  input [18:0] Wgt_3_645, // sfix19_En18
  input [18:0] Wgt_3_646, // sfix19_En18
  input [18:0] Wgt_3_647, // sfix19_En18
  input [18:0] Wgt_3_648, // sfix19_En18
  input [18:0] Wgt_3_649, // sfix19_En18
  input [18:0] Wgt_3_650, // sfix19_En18
  input [18:0] Wgt_3_651, // sfix19_En18
  input [18:0] Wgt_3_652, // sfix19_En18
  input [18:0] Wgt_3_653, // sfix19_En18
  input [18:0] Wgt_3_654, // sfix19_En18
  input [18:0] Wgt_3_655, // sfix19_En18
  input [18:0] Wgt_3_656, // sfix19_En18
  input [18:0] Wgt_3_657, // sfix19_En18
  input [18:0] Wgt_3_658, // sfix19_En18
  input [18:0] Wgt_3_659, // sfix19_En18
  input [18:0] Wgt_3_660, // sfix19_En18
  input [18:0] Wgt_3_661, // sfix19_En18
  input [18:0] Wgt_3_662, // sfix19_En18
  input [18:0] Wgt_3_663, // sfix19_En18
  input [18:0] Wgt_3_664, // sfix19_En18
  input [18:0] Wgt_3_665, // sfix19_En18
  input [18:0] Wgt_3_666, // sfix19_En18
  input [18:0] Wgt_3_667, // sfix19_En18
  input [18:0] Wgt_3_668, // sfix19_En18
  input [18:0] Wgt_3_669, // sfix19_En18
  input [18:0] Wgt_3_670, // sfix19_En18
  input [18:0] Wgt_3_671, // sfix19_En18
  input [18:0] Wgt_3_672, // sfix19_En18
  input [18:0] Wgt_3_673, // sfix19_En18
  input [18:0] Wgt_3_674, // sfix19_En18
  input [18:0] Wgt_3_675, // sfix19_En18
  input [18:0] Wgt_3_676, // sfix19_En18
  input [18:0] Wgt_3_677, // sfix19_En18
  input [18:0] Wgt_3_678, // sfix19_En18
  input [18:0] Wgt_3_679, // sfix19_En18
  input [18:0] Wgt_3_680, // sfix19_En18
  input [18:0] Wgt_3_681, // sfix19_En18
  input [18:0] Wgt_3_682, // sfix19_En18
  input [18:0] Wgt_3_683, // sfix19_En18
  input [18:0] Wgt_3_684, // sfix19_En18
  input [18:0] Wgt_3_685, // sfix19_En18
  input [18:0] Wgt_3_686, // sfix19_En18
  input [18:0] Wgt_3_687, // sfix19_En18
  input [18:0] Wgt_3_688, // sfix19_En18
  input [18:0] Wgt_3_689, // sfix19_En18
  input [18:0] Wgt_3_690, // sfix19_En18
  input [18:0] Wgt_3_691, // sfix19_En18
  input [18:0] Wgt_3_692, // sfix19_En18
  input [18:0] Wgt_3_693, // sfix19_En18
  input [18:0] Wgt_3_694, // sfix19_En18
  input [18:0] Wgt_3_695, // sfix19_En18
  input [18:0] Wgt_3_696, // sfix19_En18
  input [18:0] Wgt_3_697, // sfix19_En18
  input [18:0] Wgt_3_698, // sfix19_En18
  input [18:0] Wgt_3_699, // sfix19_En18
  input [18:0] Wgt_3_700, // sfix19_En18
  input [18:0] Wgt_3_701, // sfix19_En18
  input [18:0] Wgt_3_702, // sfix19_En18
  input [18:0] Wgt_3_703, // sfix19_En18
  input [18:0] Wgt_3_704, // sfix19_En18
  input [18:0] Wgt_3_705, // sfix19_En18
  input [18:0] Wgt_3_706, // sfix19_En18
  input [18:0] Wgt_3_707, // sfix19_En18
  input [18:0] Wgt_3_708, // sfix19_En18
  input [18:0] Wgt_3_709, // sfix19_En18
  input [18:0] Wgt_3_710, // sfix19_En18
  input [18:0] Wgt_3_711, // sfix19_En18
  input [18:0] Wgt_3_712, // sfix19_En18
  input [18:0] Wgt_3_713, // sfix19_En18
  input [18:0] Wgt_3_714, // sfix19_En18
  input [18:0] Wgt_3_715, // sfix19_En18
  input [18:0] Wgt_3_716, // sfix19_En18
  input [18:0] Wgt_3_717, // sfix19_En18
  input [18:0] Wgt_3_718, // sfix19_En18
  input [18:0] Wgt_3_719, // sfix19_En18
  input [18:0] Wgt_3_720, // sfix19_En18
  input [18:0] Wgt_3_721, // sfix19_En18
  input [18:0] Wgt_3_722, // sfix19_En18
  input [18:0] Wgt_3_723, // sfix19_En18
  input [18:0] Wgt_3_724, // sfix19_En18
  input [18:0] Wgt_3_725, // sfix19_En18
  input [18:0] Wgt_3_726, // sfix19_En18
  input [18:0] Wgt_3_727, // sfix19_En18
  input [18:0] Wgt_3_728, // sfix19_En18
  input [18:0] Wgt_3_729, // sfix19_En18
  input [18:0] Wgt_3_730, // sfix19_En18
  input [18:0] Wgt_3_731, // sfix19_En18
  input [18:0] Wgt_3_732, // sfix19_En18
  input [18:0] Wgt_3_733, // sfix19_En18
  input [18:0] Wgt_3_734, // sfix19_En18
  input [18:0] Wgt_3_735, // sfix19_En18
  input [18:0] Wgt_3_736, // sfix19_En18
  input [18:0] Wgt_3_737, // sfix19_En18
  input [18:0] Wgt_3_738, // sfix19_En18
  input [18:0] Wgt_3_739, // sfix19_En18
  input [18:0] Wgt_3_740, // sfix19_En18
  input [18:0] Wgt_3_741, // sfix19_En18
  input [18:0] Wgt_3_742, // sfix19_En18
  input [18:0] Wgt_3_743, // sfix19_En18
  input [18:0] Wgt_3_744, // sfix19_En18
  input [18:0] Wgt_3_745, // sfix19_En18
  input [18:0] Wgt_3_746, // sfix19_En18
  input [18:0] Wgt_3_747, // sfix19_En18
  input [18:0] Wgt_3_748, // sfix19_En18
  input [18:0] Wgt_3_749, // sfix19_En18
  input [18:0] Wgt_3_750, // sfix19_En18
  input [18:0] Wgt_3_751, // sfix19_En18
  input [18:0] Wgt_3_752, // sfix19_En18
  input [18:0] Wgt_3_753, // sfix19_En18
  input [18:0] Wgt_3_754, // sfix19_En18
  input [18:0] Wgt_3_755, // sfix19_En18
  input [18:0] Wgt_3_756, // sfix19_En18
  input [18:0] Wgt_3_757, // sfix19_En18
  input [18:0] Wgt_3_758, // sfix19_En18
  input [18:0] Wgt_3_759, // sfix19_En18
  input [18:0] Wgt_3_760, // sfix19_En18
  input [18:0] Wgt_3_761, // sfix19_En18
  input [18:0] Wgt_3_762, // sfix19_En18
  input [18:0] Wgt_3_763, // sfix19_En18
  input [18:0] Wgt_3_764, // sfix19_En18
  input [18:0] Wgt_3_765, // sfix19_En18
  input [18:0] Wgt_3_766, // sfix19_En18
  input [18:0] Wgt_3_767, // sfix19_En18
  input [18:0] Wgt_3_768, // sfix19_En18
  input [18:0] Wgt_3_769, // sfix19_En18
  input [18:0] Wgt_3_770, // sfix19_En18
  input [18:0] Wgt_3_771, // sfix19_En18
  input [18:0] Wgt_3_772, // sfix19_En18
  input [18:0] Wgt_3_773, // sfix19_En18
  input [18:0] Wgt_3_774, // sfix19_En18
  input [18:0] Wgt_3_775, // sfix19_En18
  input [18:0] Wgt_3_776, // sfix19_En18
  input [18:0] Wgt_3_777, // sfix19_En18
  input [18:0] Wgt_3_778, // sfix19_En18
  input [18:0] Wgt_3_779, // sfix19_En18
  input [18:0] Wgt_3_780, // sfix19_En18
  input [18:0] Wgt_3_781, // sfix19_En18
  input [18:0] Wgt_3_782, // sfix19_En18
  input [18:0] Wgt_3_783, // sfix19_En18
  input [18:0] Wgt_3_784, // sfix19_En18
  input [18:0] Wgt_4_0, // sfix19_En18
  input [18:0] Wgt_4_1, // sfix19_En18
  input [18:0] Wgt_4_2, // sfix19_En18
  input [18:0] Wgt_4_3, // sfix19_En18
  input [18:0] Wgt_4_4, // sfix19_En18
  input [18:0] Wgt_4_5, // sfix19_En18
  input [18:0] Wgt_4_6, // sfix19_En18
  input [18:0] Wgt_4_7, // sfix19_En18
  input [18:0] Wgt_4_8, // sfix19_En18
  input [18:0] Wgt_4_9, // sfix19_En18
  input [18:0] Wgt_4_10, // sfix19_En18
  input [18:0] Wgt_4_11, // sfix19_En18
  input [18:0] Wgt_4_12, // sfix19_En18
  input [18:0] Wgt_4_13, // sfix19_En18
  input [18:0] Wgt_4_14, // sfix19_En18
  input [18:0] Wgt_4_15, // sfix19_En18
  input [18:0] Wgt_4_16, // sfix19_En18
  input [18:0] Wgt_4_17, // sfix19_En18
  input [18:0] Wgt_4_18, // sfix19_En18
  input [18:0] Wgt_4_19, // sfix19_En18
  input [18:0] Wgt_4_20, // sfix19_En18
  input [18:0] Wgt_4_21, // sfix19_En18
  input [18:0] Wgt_4_22, // sfix19_En18
  input [18:0] Wgt_4_23, // sfix19_En18
  input [18:0] Wgt_4_24, // sfix19_En18
  input [18:0] Wgt_4_25, // sfix19_En18
  input [18:0] Wgt_4_26, // sfix19_En18
  input [18:0] Wgt_4_27, // sfix19_En18
  input [18:0] Wgt_4_28, // sfix19_En18
  input [18:0] Wgt_4_29, // sfix19_En18
  input [18:0] Wgt_4_30, // sfix19_En18
  input [18:0] Wgt_4_31, // sfix19_En18
  input [18:0] Wgt_4_32, // sfix19_En18
  input [18:0] Wgt_4_33, // sfix19_En18
  input [18:0] Wgt_4_34, // sfix19_En18
  input [18:0] Wgt_4_35, // sfix19_En18
  input [18:0] Wgt_4_36, // sfix19_En18
  input [18:0] Wgt_4_37, // sfix19_En18
  input [18:0] Wgt_4_38, // sfix19_En18
  input [18:0] Wgt_4_39, // sfix19_En18
  input [18:0] Wgt_4_40, // sfix19_En18
  input [18:0] Wgt_4_41, // sfix19_En18
  input [18:0] Wgt_4_42, // sfix19_En18
  input [18:0] Wgt_4_43, // sfix19_En18
  input [18:0] Wgt_4_44, // sfix19_En18
  input [18:0] Wgt_4_45, // sfix19_En18
  input [18:0] Wgt_4_46, // sfix19_En18
  input [18:0] Wgt_4_47, // sfix19_En18
  input [18:0] Wgt_4_48, // sfix19_En18
  input [18:0] Wgt_4_49, // sfix19_En18
  input [18:0] Wgt_4_50, // sfix19_En18
  input [18:0] Wgt_4_51, // sfix19_En18
  input [18:0] Wgt_4_52, // sfix19_En18
  input [18:0] Wgt_4_53, // sfix19_En18
  input [18:0] Wgt_4_54, // sfix19_En18
  input [18:0] Wgt_4_55, // sfix19_En18
  input [18:0] Wgt_4_56, // sfix19_En18
  input [18:0] Wgt_4_57, // sfix19_En18
  input [18:0] Wgt_4_58, // sfix19_En18
  input [18:0] Wgt_4_59, // sfix19_En18
  input [18:0] Wgt_4_60, // sfix19_En18
  input [18:0] Wgt_4_61, // sfix19_En18
  input [18:0] Wgt_4_62, // sfix19_En18
  input [18:0] Wgt_4_63, // sfix19_En18
  input [18:0] Wgt_4_64, // sfix19_En18
  input [18:0] Wgt_4_65, // sfix19_En18
  input [18:0] Wgt_4_66, // sfix19_En18
  input [18:0] Wgt_4_67, // sfix19_En18
  input [18:0] Wgt_4_68, // sfix19_En18
  input [18:0] Wgt_4_69, // sfix19_En18
  input [18:0] Wgt_4_70, // sfix19_En18
  input [18:0] Wgt_4_71, // sfix19_En18
  input [18:0] Wgt_4_72, // sfix19_En18
  input [18:0] Wgt_4_73, // sfix19_En18
  input [18:0] Wgt_4_74, // sfix19_En18
  input [18:0] Wgt_4_75, // sfix19_En18
  input [18:0] Wgt_4_76, // sfix19_En18
  input [18:0] Wgt_4_77, // sfix19_En18
  input [18:0] Wgt_4_78, // sfix19_En18
  input [18:0] Wgt_4_79, // sfix19_En18
  input [18:0] Wgt_4_80, // sfix19_En18
  input [18:0] Wgt_4_81, // sfix19_En18
  input [18:0] Wgt_4_82, // sfix19_En18
  input [18:0] Wgt_4_83, // sfix19_En18
  input [18:0] Wgt_4_84, // sfix19_En18
  input [18:0] Wgt_4_85, // sfix19_En18
  input [18:0] Wgt_4_86, // sfix19_En18
  input [18:0] Wgt_4_87, // sfix19_En18
  input [18:0] Wgt_4_88, // sfix19_En18
  input [18:0] Wgt_4_89, // sfix19_En18
  input [18:0] Wgt_4_90, // sfix19_En18
  input [18:0] Wgt_4_91, // sfix19_En18
  input [18:0] Wgt_4_92, // sfix19_En18
  input [18:0] Wgt_4_93, // sfix19_En18
  input [18:0] Wgt_4_94, // sfix19_En18
  input [18:0] Wgt_4_95, // sfix19_En18
  input [18:0] Wgt_4_96, // sfix19_En18
  input [18:0] Wgt_4_97, // sfix19_En18
  input [18:0] Wgt_4_98, // sfix19_En18
  input [18:0] Wgt_4_99, // sfix19_En18
  input [18:0] Wgt_4_100, // sfix19_En18
  input [18:0] Wgt_4_101, // sfix19_En18
  input [18:0] Wgt_4_102, // sfix19_En18
  input [18:0] Wgt_4_103, // sfix19_En18
  input [18:0] Wgt_4_104, // sfix19_En18
  input [18:0] Wgt_4_105, // sfix19_En18
  input [18:0] Wgt_4_106, // sfix19_En18
  input [18:0] Wgt_4_107, // sfix19_En18
  input [18:0] Wgt_4_108, // sfix19_En18
  input [18:0] Wgt_4_109, // sfix19_En18
  input [18:0] Wgt_4_110, // sfix19_En18
  input [18:0] Wgt_4_111, // sfix19_En18
  input [18:0] Wgt_4_112, // sfix19_En18
  input [18:0] Wgt_4_113, // sfix19_En18
  input [18:0] Wgt_4_114, // sfix19_En18
  input [18:0] Wgt_4_115, // sfix19_En18
  input [18:0] Wgt_4_116, // sfix19_En18
  input [18:0] Wgt_4_117, // sfix19_En18
  input [18:0] Wgt_4_118, // sfix19_En18
  input [18:0] Wgt_4_119, // sfix19_En18
  input [18:0] Wgt_4_120, // sfix19_En18
  input [18:0] Wgt_4_121, // sfix19_En18
  input [18:0] Wgt_4_122, // sfix19_En18
  input [18:0] Wgt_4_123, // sfix19_En18
  input [18:0] Wgt_4_124, // sfix19_En18
  input [18:0] Wgt_4_125, // sfix19_En18
  input [18:0] Wgt_4_126, // sfix19_En18
  input [18:0] Wgt_4_127, // sfix19_En18
  input [18:0] Wgt_4_128, // sfix19_En18
  input [18:0] Wgt_4_129, // sfix19_En18
  input [18:0] Wgt_4_130, // sfix19_En18
  input [18:0] Wgt_4_131, // sfix19_En18
  input [18:0] Wgt_4_132, // sfix19_En18
  input [18:0] Wgt_4_133, // sfix19_En18
  input [18:0] Wgt_4_134, // sfix19_En18
  input [18:0] Wgt_4_135, // sfix19_En18
  input [18:0] Wgt_4_136, // sfix19_En18
  input [18:0] Wgt_4_137, // sfix19_En18
  input [18:0] Wgt_4_138, // sfix19_En18
  input [18:0] Wgt_4_139, // sfix19_En18
  input [18:0] Wgt_4_140, // sfix19_En18
  input [18:0] Wgt_4_141, // sfix19_En18
  input [18:0] Wgt_4_142, // sfix19_En18
  input [18:0] Wgt_4_143, // sfix19_En18
  input [18:0] Wgt_4_144, // sfix19_En18
  input [18:0] Wgt_4_145, // sfix19_En18
  input [18:0] Wgt_4_146, // sfix19_En18
  input [18:0] Wgt_4_147, // sfix19_En18
  input [18:0] Wgt_4_148, // sfix19_En18
  input [18:0] Wgt_4_149, // sfix19_En18
  input [18:0] Wgt_4_150, // sfix19_En18
  input [18:0] Wgt_4_151, // sfix19_En18
  input [18:0] Wgt_4_152, // sfix19_En18
  input [18:0] Wgt_4_153, // sfix19_En18
  input [18:0] Wgt_4_154, // sfix19_En18
  input [18:0] Wgt_4_155, // sfix19_En18
  input [18:0] Wgt_4_156, // sfix19_En18
  input [18:0] Wgt_4_157, // sfix19_En18
  input [18:0] Wgt_4_158, // sfix19_En18
  input [18:0] Wgt_4_159, // sfix19_En18
  input [18:0] Wgt_4_160, // sfix19_En18
  input [18:0] Wgt_4_161, // sfix19_En18
  input [18:0] Wgt_4_162, // sfix19_En18
  input [18:0] Wgt_4_163, // sfix19_En18
  input [18:0] Wgt_4_164, // sfix19_En18
  input [18:0] Wgt_4_165, // sfix19_En18
  input [18:0] Wgt_4_166, // sfix19_En18
  input [18:0] Wgt_4_167, // sfix19_En18
  input [18:0] Wgt_4_168, // sfix19_En18
  input [18:0] Wgt_4_169, // sfix19_En18
  input [18:0] Wgt_4_170, // sfix19_En18
  input [18:0] Wgt_4_171, // sfix19_En18
  input [18:0] Wgt_4_172, // sfix19_En18
  input [18:0] Wgt_4_173, // sfix19_En18
  input [18:0] Wgt_4_174, // sfix19_En18
  input [18:0] Wgt_4_175, // sfix19_En18
  input [18:0] Wgt_4_176, // sfix19_En18
  input [18:0] Wgt_4_177, // sfix19_En18
  input [18:0] Wgt_4_178, // sfix19_En18
  input [18:0] Wgt_4_179, // sfix19_En18
  input [18:0] Wgt_4_180, // sfix19_En18
  input [18:0] Wgt_4_181, // sfix19_En18
  input [18:0] Wgt_4_182, // sfix19_En18
  input [18:0] Wgt_4_183, // sfix19_En18
  input [18:0] Wgt_4_184, // sfix19_En18
  input [18:0] Wgt_4_185, // sfix19_En18
  input [18:0] Wgt_4_186, // sfix19_En18
  input [18:0] Wgt_4_187, // sfix19_En18
  input [18:0] Wgt_4_188, // sfix19_En18
  input [18:0] Wgt_4_189, // sfix19_En18
  input [18:0] Wgt_4_190, // sfix19_En18
  input [18:0] Wgt_4_191, // sfix19_En18
  input [18:0] Wgt_4_192, // sfix19_En18
  input [18:0] Wgt_4_193, // sfix19_En18
  input [18:0] Wgt_4_194, // sfix19_En18
  input [18:0] Wgt_4_195, // sfix19_En18
  input [18:0] Wgt_4_196, // sfix19_En18
  input [18:0] Wgt_4_197, // sfix19_En18
  input [18:0] Wgt_4_198, // sfix19_En18
  input [18:0] Wgt_4_199, // sfix19_En18
  input [18:0] Wgt_4_200, // sfix19_En18
  input [18:0] Wgt_4_201, // sfix19_En18
  input [18:0] Wgt_4_202, // sfix19_En18
  input [18:0] Wgt_4_203, // sfix19_En18
  input [18:0] Wgt_4_204, // sfix19_En18
  input [18:0] Wgt_4_205, // sfix19_En18
  input [18:0] Wgt_4_206, // sfix19_En18
  input [18:0] Wgt_4_207, // sfix19_En18
  input [18:0] Wgt_4_208, // sfix19_En18
  input [18:0] Wgt_4_209, // sfix19_En18
  input [18:0] Wgt_4_210, // sfix19_En18
  input [18:0] Wgt_4_211, // sfix19_En18
  input [18:0] Wgt_4_212, // sfix19_En18
  input [18:0] Wgt_4_213, // sfix19_En18
  input [18:0] Wgt_4_214, // sfix19_En18
  input [18:0] Wgt_4_215, // sfix19_En18
  input [18:0] Wgt_4_216, // sfix19_En18
  input [18:0] Wgt_4_217, // sfix19_En18
  input [18:0] Wgt_4_218, // sfix19_En18
  input [18:0] Wgt_4_219, // sfix19_En18
  input [18:0] Wgt_4_220, // sfix19_En18
  input [18:0] Wgt_4_221, // sfix19_En18
  input [18:0] Wgt_4_222, // sfix19_En18
  input [18:0] Wgt_4_223, // sfix19_En18
  input [18:0] Wgt_4_224, // sfix19_En18
  input [18:0] Wgt_4_225, // sfix19_En18
  input [18:0] Wgt_4_226, // sfix19_En18
  input [18:0] Wgt_4_227, // sfix19_En18
  input [18:0] Wgt_4_228, // sfix19_En18
  input [18:0] Wgt_4_229, // sfix19_En18
  input [18:0] Wgt_4_230, // sfix19_En18
  input [18:0] Wgt_4_231, // sfix19_En18
  input [18:0] Wgt_4_232, // sfix19_En18
  input [18:0] Wgt_4_233, // sfix19_En18
  input [18:0] Wgt_4_234, // sfix19_En18
  input [18:0] Wgt_4_235, // sfix19_En18
  input [18:0] Wgt_4_236, // sfix19_En18
  input [18:0] Wgt_4_237, // sfix19_En18
  input [18:0] Wgt_4_238, // sfix19_En18
  input [18:0] Wgt_4_239, // sfix19_En18
  input [18:0] Wgt_4_240, // sfix19_En18
  input [18:0] Wgt_4_241, // sfix19_En18
  input [18:0] Wgt_4_242, // sfix19_En18
  input [18:0] Wgt_4_243, // sfix19_En18
  input [18:0] Wgt_4_244, // sfix19_En18
  input [18:0] Wgt_4_245, // sfix19_En18
  input [18:0] Wgt_4_246, // sfix19_En18
  input [18:0] Wgt_4_247, // sfix19_En18
  input [18:0] Wgt_4_248, // sfix19_En18
  input [18:0] Wgt_4_249, // sfix19_En18
  input [18:0] Wgt_4_250, // sfix19_En18
  input [18:0] Wgt_4_251, // sfix19_En18
  input [18:0] Wgt_4_252, // sfix19_En18
  input [18:0] Wgt_4_253, // sfix19_En18
  input [18:0] Wgt_4_254, // sfix19_En18
  input [18:0] Wgt_4_255, // sfix19_En18
  input [18:0] Wgt_4_256, // sfix19_En18
  input [18:0] Wgt_4_257, // sfix19_En18
  input [18:0] Wgt_4_258, // sfix19_En18
  input [18:0] Wgt_4_259, // sfix19_En18
  input [18:0] Wgt_4_260, // sfix19_En18
  input [18:0] Wgt_4_261, // sfix19_En18
  input [18:0] Wgt_4_262, // sfix19_En18
  input [18:0] Wgt_4_263, // sfix19_En18
  input [18:0] Wgt_4_264, // sfix19_En18
  input [18:0] Wgt_4_265, // sfix19_En18
  input [18:0] Wgt_4_266, // sfix19_En18
  input [18:0] Wgt_4_267, // sfix19_En18
  input [18:0] Wgt_4_268, // sfix19_En18
  input [18:0] Wgt_4_269, // sfix19_En18
  input [18:0] Wgt_4_270, // sfix19_En18
  input [18:0] Wgt_4_271, // sfix19_En18
  input [18:0] Wgt_4_272, // sfix19_En18
  input [18:0] Wgt_4_273, // sfix19_En18
  input [18:0] Wgt_4_274, // sfix19_En18
  input [18:0] Wgt_4_275, // sfix19_En18
  input [18:0] Wgt_4_276, // sfix19_En18
  input [18:0] Wgt_4_277, // sfix19_En18
  input [18:0] Wgt_4_278, // sfix19_En18
  input [18:0] Wgt_4_279, // sfix19_En18
  input [18:0] Wgt_4_280, // sfix19_En18
  input [18:0] Wgt_4_281, // sfix19_En18
  input [18:0] Wgt_4_282, // sfix19_En18
  input [18:0] Wgt_4_283, // sfix19_En18
  input [18:0] Wgt_4_284, // sfix19_En18
  input [18:0] Wgt_4_285, // sfix19_En18
  input [18:0] Wgt_4_286, // sfix19_En18
  input [18:0] Wgt_4_287, // sfix19_En18
  input [18:0] Wgt_4_288, // sfix19_En18
  input [18:0] Wgt_4_289, // sfix19_En18
  input [18:0] Wgt_4_290, // sfix19_En18
  input [18:0] Wgt_4_291, // sfix19_En18
  input [18:0] Wgt_4_292, // sfix19_En18
  input [18:0] Wgt_4_293, // sfix19_En18
  input [18:0] Wgt_4_294, // sfix19_En18
  input [18:0] Wgt_4_295, // sfix19_En18
  input [18:0] Wgt_4_296, // sfix19_En18
  input [18:0] Wgt_4_297, // sfix19_En18
  input [18:0] Wgt_4_298, // sfix19_En18
  input [18:0] Wgt_4_299, // sfix19_En18
  input [18:0] Wgt_4_300, // sfix19_En18
  input [18:0] Wgt_4_301, // sfix19_En18
  input [18:0] Wgt_4_302, // sfix19_En18
  input [18:0] Wgt_4_303, // sfix19_En18
  input [18:0] Wgt_4_304, // sfix19_En18
  input [18:0] Wgt_4_305, // sfix19_En18
  input [18:0] Wgt_4_306, // sfix19_En18
  input [18:0] Wgt_4_307, // sfix19_En18
  input [18:0] Wgt_4_308, // sfix19_En18
  input [18:0] Wgt_4_309, // sfix19_En18
  input [18:0] Wgt_4_310, // sfix19_En18
  input [18:0] Wgt_4_311, // sfix19_En18
  input [18:0] Wgt_4_312, // sfix19_En18
  input [18:0] Wgt_4_313, // sfix19_En18
  input [18:0] Wgt_4_314, // sfix19_En18
  input [18:0] Wgt_4_315, // sfix19_En18
  input [18:0] Wgt_4_316, // sfix19_En18
  input [18:0] Wgt_4_317, // sfix19_En18
  input [18:0] Wgt_4_318, // sfix19_En18
  input [18:0] Wgt_4_319, // sfix19_En18
  input [18:0] Wgt_4_320, // sfix19_En18
  input [18:0] Wgt_4_321, // sfix19_En18
  input [18:0] Wgt_4_322, // sfix19_En18
  input [18:0] Wgt_4_323, // sfix19_En18
  input [18:0] Wgt_4_324, // sfix19_En18
  input [18:0] Wgt_4_325, // sfix19_En18
  input [18:0] Wgt_4_326, // sfix19_En18
  input [18:0] Wgt_4_327, // sfix19_En18
  input [18:0] Wgt_4_328, // sfix19_En18
  input [18:0] Wgt_4_329, // sfix19_En18
  input [18:0] Wgt_4_330, // sfix19_En18
  input [18:0] Wgt_4_331, // sfix19_En18
  input [18:0] Wgt_4_332, // sfix19_En18
  input [18:0] Wgt_4_333, // sfix19_En18
  input [18:0] Wgt_4_334, // sfix19_En18
  input [18:0] Wgt_4_335, // sfix19_En18
  input [18:0] Wgt_4_336, // sfix19_En18
  input [18:0] Wgt_4_337, // sfix19_En18
  input [18:0] Wgt_4_338, // sfix19_En18
  input [18:0] Wgt_4_339, // sfix19_En18
  input [18:0] Wgt_4_340, // sfix19_En18
  input [18:0] Wgt_4_341, // sfix19_En18
  input [18:0] Wgt_4_342, // sfix19_En18
  input [18:0] Wgt_4_343, // sfix19_En18
  input [18:0] Wgt_4_344, // sfix19_En18
  input [18:0] Wgt_4_345, // sfix19_En18
  input [18:0] Wgt_4_346, // sfix19_En18
  input [18:0] Wgt_4_347, // sfix19_En18
  input [18:0] Wgt_4_348, // sfix19_En18
  input [18:0] Wgt_4_349, // sfix19_En18
  input [18:0] Wgt_4_350, // sfix19_En18
  input [18:0] Wgt_4_351, // sfix19_En18
  input [18:0] Wgt_4_352, // sfix19_En18
  input [18:0] Wgt_4_353, // sfix19_En18
  input [18:0] Wgt_4_354, // sfix19_En18
  input [18:0] Wgt_4_355, // sfix19_En18
  input [18:0] Wgt_4_356, // sfix19_En18
  input [18:0] Wgt_4_357, // sfix19_En18
  input [18:0] Wgt_4_358, // sfix19_En18
  input [18:0] Wgt_4_359, // sfix19_En18
  input [18:0] Wgt_4_360, // sfix19_En18
  input [18:0] Wgt_4_361, // sfix19_En18
  input [18:0] Wgt_4_362, // sfix19_En18
  input [18:0] Wgt_4_363, // sfix19_En18
  input [18:0] Wgt_4_364, // sfix19_En18
  input [18:0] Wgt_4_365, // sfix19_En18
  input [18:0] Wgt_4_366, // sfix19_En18
  input [18:0] Wgt_4_367, // sfix19_En18
  input [18:0] Wgt_4_368, // sfix19_En18
  input [18:0] Wgt_4_369, // sfix19_En18
  input [18:0] Wgt_4_370, // sfix19_En18
  input [18:0] Wgt_4_371, // sfix19_En18
  input [18:0] Wgt_4_372, // sfix19_En18
  input [18:0] Wgt_4_373, // sfix19_En18
  input [18:0] Wgt_4_374, // sfix19_En18
  input [18:0] Wgt_4_375, // sfix19_En18
  input [18:0] Wgt_4_376, // sfix19_En18
  input [18:0] Wgt_4_377, // sfix19_En18
  input [18:0] Wgt_4_378, // sfix19_En18
  input [18:0] Wgt_4_379, // sfix19_En18
  input [18:0] Wgt_4_380, // sfix19_En18
  input [18:0] Wgt_4_381, // sfix19_En18
  input [18:0] Wgt_4_382, // sfix19_En18
  input [18:0] Wgt_4_383, // sfix19_En18
  input [18:0] Wgt_4_384, // sfix19_En18
  input [18:0] Wgt_4_385, // sfix19_En18
  input [18:0] Wgt_4_386, // sfix19_En18
  input [18:0] Wgt_4_387, // sfix19_En18
  input [18:0] Wgt_4_388, // sfix19_En18
  input [18:0] Wgt_4_389, // sfix19_En18
  input [18:0] Wgt_4_390, // sfix19_En18
  input [18:0] Wgt_4_391, // sfix19_En18
  input [18:0] Wgt_4_392, // sfix19_En18
  input [18:0] Wgt_4_393, // sfix19_En18
  input [18:0] Wgt_4_394, // sfix19_En18
  input [18:0] Wgt_4_395, // sfix19_En18
  input [18:0] Wgt_4_396, // sfix19_En18
  input [18:0] Wgt_4_397, // sfix19_En18
  input [18:0] Wgt_4_398, // sfix19_En18
  input [18:0] Wgt_4_399, // sfix19_En18
  input [18:0] Wgt_4_400, // sfix19_En18
  input [18:0] Wgt_4_401, // sfix19_En18
  input [18:0] Wgt_4_402, // sfix19_En18
  input [18:0] Wgt_4_403, // sfix19_En18
  input [18:0] Wgt_4_404, // sfix19_En18
  input [18:0] Wgt_4_405, // sfix19_En18
  input [18:0] Wgt_4_406, // sfix19_En18
  input [18:0] Wgt_4_407, // sfix19_En18
  input [18:0] Wgt_4_408, // sfix19_En18
  input [18:0] Wgt_4_409, // sfix19_En18
  input [18:0] Wgt_4_410, // sfix19_En18
  input [18:0] Wgt_4_411, // sfix19_En18
  input [18:0] Wgt_4_412, // sfix19_En18
  input [18:0] Wgt_4_413, // sfix19_En18
  input [18:0] Wgt_4_414, // sfix19_En18
  input [18:0] Wgt_4_415, // sfix19_En18
  input [18:0] Wgt_4_416, // sfix19_En18
  input [18:0] Wgt_4_417, // sfix19_En18
  input [18:0] Wgt_4_418, // sfix19_En18
  input [18:0] Wgt_4_419, // sfix19_En18
  input [18:0] Wgt_4_420, // sfix19_En18
  input [18:0] Wgt_4_421, // sfix19_En18
  input [18:0] Wgt_4_422, // sfix19_En18
  input [18:0] Wgt_4_423, // sfix19_En18
  input [18:0] Wgt_4_424, // sfix19_En18
  input [18:0] Wgt_4_425, // sfix19_En18
  input [18:0] Wgt_4_426, // sfix19_En18
  input [18:0] Wgt_4_427, // sfix19_En18
  input [18:0] Wgt_4_428, // sfix19_En18
  input [18:0] Wgt_4_429, // sfix19_En18
  input [18:0] Wgt_4_430, // sfix19_En18
  input [18:0] Wgt_4_431, // sfix19_En18
  input [18:0] Wgt_4_432, // sfix19_En18
  input [18:0] Wgt_4_433, // sfix19_En18
  input [18:0] Wgt_4_434, // sfix19_En18
  input [18:0] Wgt_4_435, // sfix19_En18
  input [18:0] Wgt_4_436, // sfix19_En18
  input [18:0] Wgt_4_437, // sfix19_En18
  input [18:0] Wgt_4_438, // sfix19_En18
  input [18:0] Wgt_4_439, // sfix19_En18
  input [18:0] Wgt_4_440, // sfix19_En18
  input [18:0] Wgt_4_441, // sfix19_En18
  input [18:0] Wgt_4_442, // sfix19_En18
  input [18:0] Wgt_4_443, // sfix19_En18
  input [18:0] Wgt_4_444, // sfix19_En18
  input [18:0] Wgt_4_445, // sfix19_En18
  input [18:0] Wgt_4_446, // sfix19_En18
  input [18:0] Wgt_4_447, // sfix19_En18
  input [18:0] Wgt_4_448, // sfix19_En18
  input [18:0] Wgt_4_449, // sfix19_En18
  input [18:0] Wgt_4_450, // sfix19_En18
  input [18:0] Wgt_4_451, // sfix19_En18
  input [18:0] Wgt_4_452, // sfix19_En18
  input [18:0] Wgt_4_453, // sfix19_En18
  input [18:0] Wgt_4_454, // sfix19_En18
  input [18:0] Wgt_4_455, // sfix19_En18
  input [18:0] Wgt_4_456, // sfix19_En18
  input [18:0] Wgt_4_457, // sfix19_En18
  input [18:0] Wgt_4_458, // sfix19_En18
  input [18:0] Wgt_4_459, // sfix19_En18
  input [18:0] Wgt_4_460, // sfix19_En18
  input [18:0] Wgt_4_461, // sfix19_En18
  input [18:0] Wgt_4_462, // sfix19_En18
  input [18:0] Wgt_4_463, // sfix19_En18
  input [18:0] Wgt_4_464, // sfix19_En18
  input [18:0] Wgt_4_465, // sfix19_En18
  input [18:0] Wgt_4_466, // sfix19_En18
  input [18:0] Wgt_4_467, // sfix19_En18
  input [18:0] Wgt_4_468, // sfix19_En18
  input [18:0] Wgt_4_469, // sfix19_En18
  input [18:0] Wgt_4_470, // sfix19_En18
  input [18:0] Wgt_4_471, // sfix19_En18
  input [18:0] Wgt_4_472, // sfix19_En18
  input [18:0] Wgt_4_473, // sfix19_En18
  input [18:0] Wgt_4_474, // sfix19_En18
  input [18:0] Wgt_4_475, // sfix19_En18
  input [18:0] Wgt_4_476, // sfix19_En18
  input [18:0] Wgt_4_477, // sfix19_En18
  input [18:0] Wgt_4_478, // sfix19_En18
  input [18:0] Wgt_4_479, // sfix19_En18
  input [18:0] Wgt_4_480, // sfix19_En18
  input [18:0] Wgt_4_481, // sfix19_En18
  input [18:0] Wgt_4_482, // sfix19_En18
  input [18:0] Wgt_4_483, // sfix19_En18
  input [18:0] Wgt_4_484, // sfix19_En18
  input [18:0] Wgt_4_485, // sfix19_En18
  input [18:0] Wgt_4_486, // sfix19_En18
  input [18:0] Wgt_4_487, // sfix19_En18
  input [18:0] Wgt_4_488, // sfix19_En18
  input [18:0] Wgt_4_489, // sfix19_En18
  input [18:0] Wgt_4_490, // sfix19_En18
  input [18:0] Wgt_4_491, // sfix19_En18
  input [18:0] Wgt_4_492, // sfix19_En18
  input [18:0] Wgt_4_493, // sfix19_En18
  input [18:0] Wgt_4_494, // sfix19_En18
  input [18:0] Wgt_4_495, // sfix19_En18
  input [18:0] Wgt_4_496, // sfix19_En18
  input [18:0] Wgt_4_497, // sfix19_En18
  input [18:0] Wgt_4_498, // sfix19_En18
  input [18:0] Wgt_4_499, // sfix19_En18
  input [18:0] Wgt_4_500, // sfix19_En18
  input [18:0] Wgt_4_501, // sfix19_En18
  input [18:0] Wgt_4_502, // sfix19_En18
  input [18:0] Wgt_4_503, // sfix19_En18
  input [18:0] Wgt_4_504, // sfix19_En18
  input [18:0] Wgt_4_505, // sfix19_En18
  input [18:0] Wgt_4_506, // sfix19_En18
  input [18:0] Wgt_4_507, // sfix19_En18
  input [18:0] Wgt_4_508, // sfix19_En18
  input [18:0] Wgt_4_509, // sfix19_En18
  input [18:0] Wgt_4_510, // sfix19_En18
  input [18:0] Wgt_4_511, // sfix19_En18
  input [18:0] Wgt_4_512, // sfix19_En18
  input [18:0] Wgt_4_513, // sfix19_En18
  input [18:0] Wgt_4_514, // sfix19_En18
  input [18:0] Wgt_4_515, // sfix19_En18
  input [18:0] Wgt_4_516, // sfix19_En18
  input [18:0] Wgt_4_517, // sfix19_En18
  input [18:0] Wgt_4_518, // sfix19_En18
  input [18:0] Wgt_4_519, // sfix19_En18
  input [18:0] Wgt_4_520, // sfix19_En18
  input [18:0] Wgt_4_521, // sfix19_En18
  input [18:0] Wgt_4_522, // sfix19_En18
  input [18:0] Wgt_4_523, // sfix19_En18
  input [18:0] Wgt_4_524, // sfix19_En18
  input [18:0] Wgt_4_525, // sfix19_En18
  input [18:0] Wgt_4_526, // sfix19_En18
  input [18:0] Wgt_4_527, // sfix19_En18
  input [18:0] Wgt_4_528, // sfix19_En18
  input [18:0] Wgt_4_529, // sfix19_En18
  input [18:0] Wgt_4_530, // sfix19_En18
  input [18:0] Wgt_4_531, // sfix19_En18
  input [18:0] Wgt_4_532, // sfix19_En18
  input [18:0] Wgt_4_533, // sfix19_En18
  input [18:0] Wgt_4_534, // sfix19_En18
  input [18:0] Wgt_4_535, // sfix19_En18
  input [18:0] Wgt_4_536, // sfix19_En18
  input [18:0] Wgt_4_537, // sfix19_En18
  input [18:0] Wgt_4_538, // sfix19_En18
  input [18:0] Wgt_4_539, // sfix19_En18
  input [18:0] Wgt_4_540, // sfix19_En18
  input [18:0] Wgt_4_541, // sfix19_En18
  input [18:0] Wgt_4_542, // sfix19_En18
  input [18:0] Wgt_4_543, // sfix19_En18
  input [18:0] Wgt_4_544, // sfix19_En18
  input [18:0] Wgt_4_545, // sfix19_En18
  input [18:0] Wgt_4_546, // sfix19_En18
  input [18:0] Wgt_4_547, // sfix19_En18
  input [18:0] Wgt_4_548, // sfix19_En18
  input [18:0] Wgt_4_549, // sfix19_En18
  input [18:0] Wgt_4_550, // sfix19_En18
  input [18:0] Wgt_4_551, // sfix19_En18
  input [18:0] Wgt_4_552, // sfix19_En18
  input [18:0] Wgt_4_553, // sfix19_En18
  input [18:0] Wgt_4_554, // sfix19_En18
  input [18:0] Wgt_4_555, // sfix19_En18
  input [18:0] Wgt_4_556, // sfix19_En18
  input [18:0] Wgt_4_557, // sfix19_En18
  input [18:0] Wgt_4_558, // sfix19_En18
  input [18:0] Wgt_4_559, // sfix19_En18
  input [18:0] Wgt_4_560, // sfix19_En18
  input [18:0] Wgt_4_561, // sfix19_En18
  input [18:0] Wgt_4_562, // sfix19_En18
  input [18:0] Wgt_4_563, // sfix19_En18
  input [18:0] Wgt_4_564, // sfix19_En18
  input [18:0] Wgt_4_565, // sfix19_En18
  input [18:0] Wgt_4_566, // sfix19_En18
  input [18:0] Wgt_4_567, // sfix19_En18
  input [18:0] Wgt_4_568, // sfix19_En18
  input [18:0] Wgt_4_569, // sfix19_En18
  input [18:0] Wgt_4_570, // sfix19_En18
  input [18:0] Wgt_4_571, // sfix19_En18
  input [18:0] Wgt_4_572, // sfix19_En18
  input [18:0] Wgt_4_573, // sfix19_En18
  input [18:0] Wgt_4_574, // sfix19_En18
  input [18:0] Wgt_4_575, // sfix19_En18
  input [18:0] Wgt_4_576, // sfix19_En18
  input [18:0] Wgt_4_577, // sfix19_En18
  input [18:0] Wgt_4_578, // sfix19_En18
  input [18:0] Wgt_4_579, // sfix19_En18
  input [18:0] Wgt_4_580, // sfix19_En18
  input [18:0] Wgt_4_581, // sfix19_En18
  input [18:0] Wgt_4_582, // sfix19_En18
  input [18:0] Wgt_4_583, // sfix19_En18
  input [18:0] Wgt_4_584, // sfix19_En18
  input [18:0] Wgt_4_585, // sfix19_En18
  input [18:0] Wgt_4_586, // sfix19_En18
  input [18:0] Wgt_4_587, // sfix19_En18
  input [18:0] Wgt_4_588, // sfix19_En18
  input [18:0] Wgt_4_589, // sfix19_En18
  input [18:0] Wgt_4_590, // sfix19_En18
  input [18:0] Wgt_4_591, // sfix19_En18
  input [18:0] Wgt_4_592, // sfix19_En18
  input [18:0] Wgt_4_593, // sfix19_En18
  input [18:0] Wgt_4_594, // sfix19_En18
  input [18:0] Wgt_4_595, // sfix19_En18
  input [18:0] Wgt_4_596, // sfix19_En18
  input [18:0] Wgt_4_597, // sfix19_En18
  input [18:0] Wgt_4_598, // sfix19_En18
  input [18:0] Wgt_4_599, // sfix19_En18
  input [18:0] Wgt_4_600, // sfix19_En18
  input [18:0] Wgt_4_601, // sfix19_En18
  input [18:0] Wgt_4_602, // sfix19_En18
  input [18:0] Wgt_4_603, // sfix19_En18
  input [18:0] Wgt_4_604, // sfix19_En18
  input [18:0] Wgt_4_605, // sfix19_En18
  input [18:0] Wgt_4_606, // sfix19_En18
  input [18:0] Wgt_4_607, // sfix19_En18
  input [18:0] Wgt_4_608, // sfix19_En18
  input [18:0] Wgt_4_609, // sfix19_En18
  input [18:0] Wgt_4_610, // sfix19_En18
  input [18:0] Wgt_4_611, // sfix19_En18
  input [18:0] Wgt_4_612, // sfix19_En18
  input [18:0] Wgt_4_613, // sfix19_En18
  input [18:0] Wgt_4_614, // sfix19_En18
  input [18:0] Wgt_4_615, // sfix19_En18
  input [18:0] Wgt_4_616, // sfix19_En18
  input [18:0] Wgt_4_617, // sfix19_En18
  input [18:0] Wgt_4_618, // sfix19_En18
  input [18:0] Wgt_4_619, // sfix19_En18
  input [18:0] Wgt_4_620, // sfix19_En18
  input [18:0] Wgt_4_621, // sfix19_En18
  input [18:0] Wgt_4_622, // sfix19_En18
  input [18:0] Wgt_4_623, // sfix19_En18
  input [18:0] Wgt_4_624, // sfix19_En18
  input [18:0] Wgt_4_625, // sfix19_En18
  input [18:0] Wgt_4_626, // sfix19_En18
  input [18:0] Wgt_4_627, // sfix19_En18
  input [18:0] Wgt_4_628, // sfix19_En18
  input [18:0] Wgt_4_629, // sfix19_En18
  input [18:0] Wgt_4_630, // sfix19_En18
  input [18:0] Wgt_4_631, // sfix19_En18
  input [18:0] Wgt_4_632, // sfix19_En18
  input [18:0] Wgt_4_633, // sfix19_En18
  input [18:0] Wgt_4_634, // sfix19_En18
  input [18:0] Wgt_4_635, // sfix19_En18
  input [18:0] Wgt_4_636, // sfix19_En18
  input [18:0] Wgt_4_637, // sfix19_En18
  input [18:0] Wgt_4_638, // sfix19_En18
  input [18:0] Wgt_4_639, // sfix19_En18
  input [18:0] Wgt_4_640, // sfix19_En18
  input [18:0] Wgt_4_641, // sfix19_En18
  input [18:0] Wgt_4_642, // sfix19_En18
  input [18:0] Wgt_4_643, // sfix19_En18
  input [18:0] Wgt_4_644, // sfix19_En18
  input [18:0] Wgt_4_645, // sfix19_En18
  input [18:0] Wgt_4_646, // sfix19_En18
  input [18:0] Wgt_4_647, // sfix19_En18
  input [18:0] Wgt_4_648, // sfix19_En18
  input [18:0] Wgt_4_649, // sfix19_En18
  input [18:0] Wgt_4_650, // sfix19_En18
  input [18:0] Wgt_4_651, // sfix19_En18
  input [18:0] Wgt_4_652, // sfix19_En18
  input [18:0] Wgt_4_653, // sfix19_En18
  input [18:0] Wgt_4_654, // sfix19_En18
  input [18:0] Wgt_4_655, // sfix19_En18
  input [18:0] Wgt_4_656, // sfix19_En18
  input [18:0] Wgt_4_657, // sfix19_En18
  input [18:0] Wgt_4_658, // sfix19_En18
  input [18:0] Wgt_4_659, // sfix19_En18
  input [18:0] Wgt_4_660, // sfix19_En18
  input [18:0] Wgt_4_661, // sfix19_En18
  input [18:0] Wgt_4_662, // sfix19_En18
  input [18:0] Wgt_4_663, // sfix19_En18
  input [18:0] Wgt_4_664, // sfix19_En18
  input [18:0] Wgt_4_665, // sfix19_En18
  input [18:0] Wgt_4_666, // sfix19_En18
  input [18:0] Wgt_4_667, // sfix19_En18
  input [18:0] Wgt_4_668, // sfix19_En18
  input [18:0] Wgt_4_669, // sfix19_En18
  input [18:0] Wgt_4_670, // sfix19_En18
  input [18:0] Wgt_4_671, // sfix19_En18
  input [18:0] Wgt_4_672, // sfix19_En18
  input [18:0] Wgt_4_673, // sfix19_En18
  input [18:0] Wgt_4_674, // sfix19_En18
  input [18:0] Wgt_4_675, // sfix19_En18
  input [18:0] Wgt_4_676, // sfix19_En18
  input [18:0] Wgt_4_677, // sfix19_En18
  input [18:0] Wgt_4_678, // sfix19_En18
  input [18:0] Wgt_4_679, // sfix19_En18
  input [18:0] Wgt_4_680, // sfix19_En18
  input [18:0] Wgt_4_681, // sfix19_En18
  input [18:0] Wgt_4_682, // sfix19_En18
  input [18:0] Wgt_4_683, // sfix19_En18
  input [18:0] Wgt_4_684, // sfix19_En18
  input [18:0] Wgt_4_685, // sfix19_En18
  input [18:0] Wgt_4_686, // sfix19_En18
  input [18:0] Wgt_4_687, // sfix19_En18
  input [18:0] Wgt_4_688, // sfix19_En18
  input [18:0] Wgt_4_689, // sfix19_En18
  input [18:0] Wgt_4_690, // sfix19_En18
  input [18:0] Wgt_4_691, // sfix19_En18
  input [18:0] Wgt_4_692, // sfix19_En18
  input [18:0] Wgt_4_693, // sfix19_En18
  input [18:0] Wgt_4_694, // sfix19_En18
  input [18:0] Wgt_4_695, // sfix19_En18
  input [18:0] Wgt_4_696, // sfix19_En18
  input [18:0] Wgt_4_697, // sfix19_En18
  input [18:0] Wgt_4_698, // sfix19_En18
  input [18:0] Wgt_4_699, // sfix19_En18
  input [18:0] Wgt_4_700, // sfix19_En18
  input [18:0] Wgt_4_701, // sfix19_En18
  input [18:0] Wgt_4_702, // sfix19_En18
  input [18:0] Wgt_4_703, // sfix19_En18
  input [18:0] Wgt_4_704, // sfix19_En18
  input [18:0] Wgt_4_705, // sfix19_En18
  input [18:0] Wgt_4_706, // sfix19_En18
  input [18:0] Wgt_4_707, // sfix19_En18
  input [18:0] Wgt_4_708, // sfix19_En18
  input [18:0] Wgt_4_709, // sfix19_En18
  input [18:0] Wgt_4_710, // sfix19_En18
  input [18:0] Wgt_4_711, // sfix19_En18
  input [18:0] Wgt_4_712, // sfix19_En18
  input [18:0] Wgt_4_713, // sfix19_En18
  input [18:0] Wgt_4_714, // sfix19_En18
  input [18:0] Wgt_4_715, // sfix19_En18
  input [18:0] Wgt_4_716, // sfix19_En18
  input [18:0] Wgt_4_717, // sfix19_En18
  input [18:0] Wgt_4_718, // sfix19_En18
  input [18:0] Wgt_4_719, // sfix19_En18
  input [18:0] Wgt_4_720, // sfix19_En18
  input [18:0] Wgt_4_721, // sfix19_En18
  input [18:0] Wgt_4_722, // sfix19_En18
  input [18:0] Wgt_4_723, // sfix19_En18
  input [18:0] Wgt_4_724, // sfix19_En18
  input [18:0] Wgt_4_725, // sfix19_En18
  input [18:0] Wgt_4_726, // sfix19_En18
  input [18:0] Wgt_4_727, // sfix19_En18
  input [18:0] Wgt_4_728, // sfix19_En18
  input [18:0] Wgt_4_729, // sfix19_En18
  input [18:0] Wgt_4_730, // sfix19_En18
  input [18:0] Wgt_4_731, // sfix19_En18
  input [18:0] Wgt_4_732, // sfix19_En18
  input [18:0] Wgt_4_733, // sfix19_En18
  input [18:0] Wgt_4_734, // sfix19_En18
  input [18:0] Wgt_4_735, // sfix19_En18
  input [18:0] Wgt_4_736, // sfix19_En18
  input [18:0] Wgt_4_737, // sfix19_En18
  input [18:0] Wgt_4_738, // sfix19_En18
  input [18:0] Wgt_4_739, // sfix19_En18
  input [18:0] Wgt_4_740, // sfix19_En18
  input [18:0] Wgt_4_741, // sfix19_En18
  input [18:0] Wgt_4_742, // sfix19_En18
  input [18:0] Wgt_4_743, // sfix19_En18
  input [18:0] Wgt_4_744, // sfix19_En18
  input [18:0] Wgt_4_745, // sfix19_En18
  input [18:0] Wgt_4_746, // sfix19_En18
  input [18:0] Wgt_4_747, // sfix19_En18
  input [18:0] Wgt_4_748, // sfix19_En18
  input [18:0] Wgt_4_749, // sfix19_En18
  input [18:0] Wgt_4_750, // sfix19_En18
  input [18:0] Wgt_4_751, // sfix19_En18
  input [18:0] Wgt_4_752, // sfix19_En18
  input [18:0] Wgt_4_753, // sfix19_En18
  input [18:0] Wgt_4_754, // sfix19_En18
  input [18:0] Wgt_4_755, // sfix19_En18
  input [18:0] Wgt_4_756, // sfix19_En18
  input [18:0] Wgt_4_757, // sfix19_En18
  input [18:0] Wgt_4_758, // sfix19_En18
  input [18:0] Wgt_4_759, // sfix19_En18
  input [18:0] Wgt_4_760, // sfix19_En18
  input [18:0] Wgt_4_761, // sfix19_En18
  input [18:0] Wgt_4_762, // sfix19_En18
  input [18:0] Wgt_4_763, // sfix19_En18
  input [18:0] Wgt_4_764, // sfix19_En18
  input [18:0] Wgt_4_765, // sfix19_En18
  input [18:0] Wgt_4_766, // sfix19_En18
  input [18:0] Wgt_4_767, // sfix19_En18
  input [18:0] Wgt_4_768, // sfix19_En18
  input [18:0] Wgt_4_769, // sfix19_En18
  input [18:0] Wgt_4_770, // sfix19_En18
  input [18:0] Wgt_4_771, // sfix19_En18
  input [18:0] Wgt_4_772, // sfix19_En18
  input [18:0] Wgt_4_773, // sfix19_En18
  input [18:0] Wgt_4_774, // sfix19_En18
  input [18:0] Wgt_4_775, // sfix19_En18
  input [18:0] Wgt_4_776, // sfix19_En18
  input [18:0] Wgt_4_777, // sfix19_En18
  input [18:0] Wgt_4_778, // sfix19_En18
  input [18:0] Wgt_4_779, // sfix19_En18
  input [18:0] Wgt_4_780, // sfix19_En18
  input [18:0] Wgt_4_781, // sfix19_En18
  input [18:0] Wgt_4_782, // sfix19_En18
  input [18:0] Wgt_4_783, // sfix19_En18
  input [18:0] Wgt_4_784, // sfix19_En18
  input [18:0] Wgt_5_0, // sfix19_En18
  input [18:0] Wgt_5_1, // sfix19_En18
  input [18:0] Wgt_5_2, // sfix19_En18
  input [18:0] Wgt_5_3, // sfix19_En18
  input [18:0] Wgt_5_4, // sfix19_En18
  input [18:0] Wgt_5_5, // sfix19_En18
  input [18:0] Wgt_5_6, // sfix19_En18
  input [18:0] Wgt_5_7, // sfix19_En18
  input [18:0] Wgt_5_8, // sfix19_En18
  input [18:0] Wgt_5_9, // sfix19_En18
  input [18:0] Wgt_5_10, // sfix19_En18
  input [18:0] Wgt_5_11, // sfix19_En18
  input [18:0] Wgt_5_12, // sfix19_En18
  input [18:0] Wgt_5_13, // sfix19_En18
  input [18:0] Wgt_5_14, // sfix19_En18
  input [18:0] Wgt_5_15, // sfix19_En18
  input [18:0] Wgt_5_16, // sfix19_En18
  input [18:0] Wgt_5_17, // sfix19_En18
  input [18:0] Wgt_5_18, // sfix19_En18
  input [18:0] Wgt_5_19, // sfix19_En18
  input [18:0] Wgt_5_20, // sfix19_En18
  input [18:0] Wgt_5_21, // sfix19_En18
  input [18:0] Wgt_5_22, // sfix19_En18
  input [18:0] Wgt_5_23, // sfix19_En18
  input [18:0] Wgt_5_24, // sfix19_En18
  input [18:0] Wgt_5_25, // sfix19_En18
  input [18:0] Wgt_5_26, // sfix19_En18
  input [18:0] Wgt_5_27, // sfix19_En18
  input [18:0] Wgt_5_28, // sfix19_En18
  input [18:0] Wgt_5_29, // sfix19_En18
  input [18:0] Wgt_5_30, // sfix19_En18
  input [18:0] Wgt_5_31, // sfix19_En18
  input [18:0] Wgt_5_32, // sfix19_En18
  input [18:0] Wgt_5_33, // sfix19_En18
  input [18:0] Wgt_5_34, // sfix19_En18
  input [18:0] Wgt_5_35, // sfix19_En18
  input [18:0] Wgt_5_36, // sfix19_En18
  input [18:0] Wgt_5_37, // sfix19_En18
  input [18:0] Wgt_5_38, // sfix19_En18
  input [18:0] Wgt_5_39, // sfix19_En18
  input [18:0] Wgt_5_40, // sfix19_En18
  input [18:0] Wgt_5_41, // sfix19_En18
  input [18:0] Wgt_5_42, // sfix19_En18
  input [18:0] Wgt_5_43, // sfix19_En18
  input [18:0] Wgt_5_44, // sfix19_En18
  input [18:0] Wgt_5_45, // sfix19_En18
  input [18:0] Wgt_5_46, // sfix19_En18
  input [18:0] Wgt_5_47, // sfix19_En18
  input [18:0] Wgt_5_48, // sfix19_En18
  input [18:0] Wgt_5_49, // sfix19_En18
  input [18:0] Wgt_5_50, // sfix19_En18
  input [18:0] Wgt_5_51, // sfix19_En18
  input [18:0] Wgt_5_52, // sfix19_En18
  input [18:0] Wgt_5_53, // sfix19_En18
  input [18:0] Wgt_5_54, // sfix19_En18
  input [18:0] Wgt_5_55, // sfix19_En18
  input [18:0] Wgt_5_56, // sfix19_En18
  input [18:0] Wgt_5_57, // sfix19_En18
  input [18:0] Wgt_5_58, // sfix19_En18
  input [18:0] Wgt_5_59, // sfix19_En18
  input [18:0] Wgt_5_60, // sfix19_En18
  input [18:0] Wgt_5_61, // sfix19_En18
  input [18:0] Wgt_5_62, // sfix19_En18
  input [18:0] Wgt_5_63, // sfix19_En18
  input [18:0] Wgt_5_64, // sfix19_En18
  input [18:0] Wgt_5_65, // sfix19_En18
  input [18:0] Wgt_5_66, // sfix19_En18
  input [18:0] Wgt_5_67, // sfix19_En18
  input [18:0] Wgt_5_68, // sfix19_En18
  input [18:0] Wgt_5_69, // sfix19_En18
  input [18:0] Wgt_5_70, // sfix19_En18
  input [18:0] Wgt_5_71, // sfix19_En18
  input [18:0] Wgt_5_72, // sfix19_En18
  input [18:0] Wgt_5_73, // sfix19_En18
  input [18:0] Wgt_5_74, // sfix19_En18
  input [18:0] Wgt_5_75, // sfix19_En18
  input [18:0] Wgt_5_76, // sfix19_En18
  input [18:0] Wgt_5_77, // sfix19_En18
  input [18:0] Wgt_5_78, // sfix19_En18
  input [18:0] Wgt_5_79, // sfix19_En18
  input [18:0] Wgt_5_80, // sfix19_En18
  input [18:0] Wgt_5_81, // sfix19_En18
  input [18:0] Wgt_5_82, // sfix19_En18
  input [18:0] Wgt_5_83, // sfix19_En18
  input [18:0] Wgt_5_84, // sfix19_En18
  input [18:0] Wgt_5_85, // sfix19_En18
  input [18:0] Wgt_5_86, // sfix19_En18
  input [18:0] Wgt_5_87, // sfix19_En18
  input [18:0] Wgt_5_88, // sfix19_En18
  input [18:0] Wgt_5_89, // sfix19_En18
  input [18:0] Wgt_5_90, // sfix19_En18
  input [18:0] Wgt_5_91, // sfix19_En18
  input [18:0] Wgt_5_92, // sfix19_En18
  input [18:0] Wgt_5_93, // sfix19_En18
  input [18:0] Wgt_5_94, // sfix19_En18
  input [18:0] Wgt_5_95, // sfix19_En18
  input [18:0] Wgt_5_96, // sfix19_En18
  input [18:0] Wgt_5_97, // sfix19_En18
  input [18:0] Wgt_5_98, // sfix19_En18
  input [18:0] Wgt_5_99, // sfix19_En18
  input [18:0] Wgt_5_100, // sfix19_En18
  input [18:0] Wgt_5_101, // sfix19_En18
  input [18:0] Wgt_5_102, // sfix19_En18
  input [18:0] Wgt_5_103, // sfix19_En18
  input [18:0] Wgt_5_104, // sfix19_En18
  input [18:0] Wgt_5_105, // sfix19_En18
  input [18:0] Wgt_5_106, // sfix19_En18
  input [18:0] Wgt_5_107, // sfix19_En18
  input [18:0] Wgt_5_108, // sfix19_En18
  input [18:0] Wgt_5_109, // sfix19_En18
  input [18:0] Wgt_5_110, // sfix19_En18
  input [18:0] Wgt_5_111, // sfix19_En18
  input [18:0] Wgt_5_112, // sfix19_En18
  input [18:0] Wgt_5_113, // sfix19_En18
  input [18:0] Wgt_5_114, // sfix19_En18
  input [18:0] Wgt_5_115, // sfix19_En18
  input [18:0] Wgt_5_116, // sfix19_En18
  input [18:0] Wgt_5_117, // sfix19_En18
  input [18:0] Wgt_5_118, // sfix19_En18
  input [18:0] Wgt_5_119, // sfix19_En18
  input [18:0] Wgt_5_120, // sfix19_En18
  input [18:0] Wgt_5_121, // sfix19_En18
  input [18:0] Wgt_5_122, // sfix19_En18
  input [18:0] Wgt_5_123, // sfix19_En18
  input [18:0] Wgt_5_124, // sfix19_En18
  input [18:0] Wgt_5_125, // sfix19_En18
  input [18:0] Wgt_5_126, // sfix19_En18
  input [18:0] Wgt_5_127, // sfix19_En18
  input [18:0] Wgt_5_128, // sfix19_En18
  input [18:0] Wgt_5_129, // sfix19_En18
  input [18:0] Wgt_5_130, // sfix19_En18
  input [18:0] Wgt_5_131, // sfix19_En18
  input [18:0] Wgt_5_132, // sfix19_En18
  input [18:0] Wgt_5_133, // sfix19_En18
  input [18:0] Wgt_5_134, // sfix19_En18
  input [18:0] Wgt_5_135, // sfix19_En18
  input [18:0] Wgt_5_136, // sfix19_En18
  input [18:0] Wgt_5_137, // sfix19_En18
  input [18:0] Wgt_5_138, // sfix19_En18
  input [18:0] Wgt_5_139, // sfix19_En18
  input [18:0] Wgt_5_140, // sfix19_En18
  input [18:0] Wgt_5_141, // sfix19_En18
  input [18:0] Wgt_5_142, // sfix19_En18
  input [18:0] Wgt_5_143, // sfix19_En18
  input [18:0] Wgt_5_144, // sfix19_En18
  input [18:0] Wgt_5_145, // sfix19_En18
  input [18:0] Wgt_5_146, // sfix19_En18
  input [18:0] Wgt_5_147, // sfix19_En18
  input [18:0] Wgt_5_148, // sfix19_En18
  input [18:0] Wgt_5_149, // sfix19_En18
  input [18:0] Wgt_5_150, // sfix19_En18
  input [18:0] Wgt_5_151, // sfix19_En18
  input [18:0] Wgt_5_152, // sfix19_En18
  input [18:0] Wgt_5_153, // sfix19_En18
  input [18:0] Wgt_5_154, // sfix19_En18
  input [18:0] Wgt_5_155, // sfix19_En18
  input [18:0] Wgt_5_156, // sfix19_En18
  input [18:0] Wgt_5_157, // sfix19_En18
  input [18:0] Wgt_5_158, // sfix19_En18
  input [18:0] Wgt_5_159, // sfix19_En18
  input [18:0] Wgt_5_160, // sfix19_En18
  input [18:0] Wgt_5_161, // sfix19_En18
  input [18:0] Wgt_5_162, // sfix19_En18
  input [18:0] Wgt_5_163, // sfix19_En18
  input [18:0] Wgt_5_164, // sfix19_En18
  input [18:0] Wgt_5_165, // sfix19_En18
  input [18:0] Wgt_5_166, // sfix19_En18
  input [18:0] Wgt_5_167, // sfix19_En18
  input [18:0] Wgt_5_168, // sfix19_En18
  input [18:0] Wgt_5_169, // sfix19_En18
  input [18:0] Wgt_5_170, // sfix19_En18
  input [18:0] Wgt_5_171, // sfix19_En18
  input [18:0] Wgt_5_172, // sfix19_En18
  input [18:0] Wgt_5_173, // sfix19_En18
  input [18:0] Wgt_5_174, // sfix19_En18
  input [18:0] Wgt_5_175, // sfix19_En18
  input [18:0] Wgt_5_176, // sfix19_En18
  input [18:0] Wgt_5_177, // sfix19_En18
  input [18:0] Wgt_5_178, // sfix19_En18
  input [18:0] Wgt_5_179, // sfix19_En18
  input [18:0] Wgt_5_180, // sfix19_En18
  input [18:0] Wgt_5_181, // sfix19_En18
  input [18:0] Wgt_5_182, // sfix19_En18
  input [18:0] Wgt_5_183, // sfix19_En18
  input [18:0] Wgt_5_184, // sfix19_En18
  input [18:0] Wgt_5_185, // sfix19_En18
  input [18:0] Wgt_5_186, // sfix19_En18
  input [18:0] Wgt_5_187, // sfix19_En18
  input [18:0] Wgt_5_188, // sfix19_En18
  input [18:0] Wgt_5_189, // sfix19_En18
  input [18:0] Wgt_5_190, // sfix19_En18
  input [18:0] Wgt_5_191, // sfix19_En18
  input [18:0] Wgt_5_192, // sfix19_En18
  input [18:0] Wgt_5_193, // sfix19_En18
  input [18:0] Wgt_5_194, // sfix19_En18
  input [18:0] Wgt_5_195, // sfix19_En18
  input [18:0] Wgt_5_196, // sfix19_En18
  input [18:0] Wgt_5_197, // sfix19_En18
  input [18:0] Wgt_5_198, // sfix19_En18
  input [18:0] Wgt_5_199, // sfix19_En18
  input [18:0] Wgt_5_200, // sfix19_En18
  input [18:0] Wgt_5_201, // sfix19_En18
  input [18:0] Wgt_5_202, // sfix19_En18
  input [18:0] Wgt_5_203, // sfix19_En18
  input [18:0] Wgt_5_204, // sfix19_En18
  input [18:0] Wgt_5_205, // sfix19_En18
  input [18:0] Wgt_5_206, // sfix19_En18
  input [18:0] Wgt_5_207, // sfix19_En18
  input [18:0] Wgt_5_208, // sfix19_En18
  input [18:0] Wgt_5_209, // sfix19_En18
  input [18:0] Wgt_5_210, // sfix19_En18
  input [18:0] Wgt_5_211, // sfix19_En18
  input [18:0] Wgt_5_212, // sfix19_En18
  input [18:0] Wgt_5_213, // sfix19_En18
  input [18:0] Wgt_5_214, // sfix19_En18
  input [18:0] Wgt_5_215, // sfix19_En18
  input [18:0] Wgt_5_216, // sfix19_En18
  input [18:0] Wgt_5_217, // sfix19_En18
  input [18:0] Wgt_5_218, // sfix19_En18
  input [18:0] Wgt_5_219, // sfix19_En18
  input [18:0] Wgt_5_220, // sfix19_En18
  input [18:0] Wgt_5_221, // sfix19_En18
  input [18:0] Wgt_5_222, // sfix19_En18
  input [18:0] Wgt_5_223, // sfix19_En18
  input [18:0] Wgt_5_224, // sfix19_En18
  input [18:0] Wgt_5_225, // sfix19_En18
  input [18:0] Wgt_5_226, // sfix19_En18
  input [18:0] Wgt_5_227, // sfix19_En18
  input [18:0] Wgt_5_228, // sfix19_En18
  input [18:0] Wgt_5_229, // sfix19_En18
  input [18:0] Wgt_5_230, // sfix19_En18
  input [18:0] Wgt_5_231, // sfix19_En18
  input [18:0] Wgt_5_232, // sfix19_En18
  input [18:0] Wgt_5_233, // sfix19_En18
  input [18:0] Wgt_5_234, // sfix19_En18
  input [18:0] Wgt_5_235, // sfix19_En18
  input [18:0] Wgt_5_236, // sfix19_En18
  input [18:0] Wgt_5_237, // sfix19_En18
  input [18:0] Wgt_5_238, // sfix19_En18
  input [18:0] Wgt_5_239, // sfix19_En18
  input [18:0] Wgt_5_240, // sfix19_En18
  input [18:0] Wgt_5_241, // sfix19_En18
  input [18:0] Wgt_5_242, // sfix19_En18
  input [18:0] Wgt_5_243, // sfix19_En18
  input [18:0] Wgt_5_244, // sfix19_En18
  input [18:0] Wgt_5_245, // sfix19_En18
  input [18:0] Wgt_5_246, // sfix19_En18
  input [18:0] Wgt_5_247, // sfix19_En18
  input [18:0] Wgt_5_248, // sfix19_En18
  input [18:0] Wgt_5_249, // sfix19_En18
  input [18:0] Wgt_5_250, // sfix19_En18
  input [18:0] Wgt_5_251, // sfix19_En18
  input [18:0] Wgt_5_252, // sfix19_En18
  input [18:0] Wgt_5_253, // sfix19_En18
  input [18:0] Wgt_5_254, // sfix19_En18
  input [18:0] Wgt_5_255, // sfix19_En18
  input [18:0] Wgt_5_256, // sfix19_En18
  input [18:0] Wgt_5_257, // sfix19_En18
  input [18:0] Wgt_5_258, // sfix19_En18
  input [18:0] Wgt_5_259, // sfix19_En18
  input [18:0] Wgt_5_260, // sfix19_En18
  input [18:0] Wgt_5_261, // sfix19_En18
  input [18:0] Wgt_5_262, // sfix19_En18
  input [18:0] Wgt_5_263, // sfix19_En18
  input [18:0] Wgt_5_264, // sfix19_En18
  input [18:0] Wgt_5_265, // sfix19_En18
  input [18:0] Wgt_5_266, // sfix19_En18
  input [18:0] Wgt_5_267, // sfix19_En18
  input [18:0] Wgt_5_268, // sfix19_En18
  input [18:0] Wgt_5_269, // sfix19_En18
  input [18:0] Wgt_5_270, // sfix19_En18
  input [18:0] Wgt_5_271, // sfix19_En18
  input [18:0] Wgt_5_272, // sfix19_En18
  input [18:0] Wgt_5_273, // sfix19_En18
  input [18:0] Wgt_5_274, // sfix19_En18
  input [18:0] Wgt_5_275, // sfix19_En18
  input [18:0] Wgt_5_276, // sfix19_En18
  input [18:0] Wgt_5_277, // sfix19_En18
  input [18:0] Wgt_5_278, // sfix19_En18
  input [18:0] Wgt_5_279, // sfix19_En18
  input [18:0] Wgt_5_280, // sfix19_En18
  input [18:0] Wgt_5_281, // sfix19_En18
  input [18:0] Wgt_5_282, // sfix19_En18
  input [18:0] Wgt_5_283, // sfix19_En18
  input [18:0] Wgt_5_284, // sfix19_En18
  input [18:0] Wgt_5_285, // sfix19_En18
  input [18:0] Wgt_5_286, // sfix19_En18
  input [18:0] Wgt_5_287, // sfix19_En18
  input [18:0] Wgt_5_288, // sfix19_En18
  input [18:0] Wgt_5_289, // sfix19_En18
  input [18:0] Wgt_5_290, // sfix19_En18
  input [18:0] Wgt_5_291, // sfix19_En18
  input [18:0] Wgt_5_292, // sfix19_En18
  input [18:0] Wgt_5_293, // sfix19_En18
  input [18:0] Wgt_5_294, // sfix19_En18
  input [18:0] Wgt_5_295, // sfix19_En18
  input [18:0] Wgt_5_296, // sfix19_En18
  input [18:0] Wgt_5_297, // sfix19_En18
  input [18:0] Wgt_5_298, // sfix19_En18
  input [18:0] Wgt_5_299, // sfix19_En18
  input [18:0] Wgt_5_300, // sfix19_En18
  input [18:0] Wgt_5_301, // sfix19_En18
  input [18:0] Wgt_5_302, // sfix19_En18
  input [18:0] Wgt_5_303, // sfix19_En18
  input [18:0] Wgt_5_304, // sfix19_En18
  input [18:0] Wgt_5_305, // sfix19_En18
  input [18:0] Wgt_5_306, // sfix19_En18
  input [18:0] Wgt_5_307, // sfix19_En18
  input [18:0] Wgt_5_308, // sfix19_En18
  input [18:0] Wgt_5_309, // sfix19_En18
  input [18:0] Wgt_5_310, // sfix19_En18
  input [18:0] Wgt_5_311, // sfix19_En18
  input [18:0] Wgt_5_312, // sfix19_En18
  input [18:0] Wgt_5_313, // sfix19_En18
  input [18:0] Wgt_5_314, // sfix19_En18
  input [18:0] Wgt_5_315, // sfix19_En18
  input [18:0] Wgt_5_316, // sfix19_En18
  input [18:0] Wgt_5_317, // sfix19_En18
  input [18:0] Wgt_5_318, // sfix19_En18
  input [18:0] Wgt_5_319, // sfix19_En18
  input [18:0] Wgt_5_320, // sfix19_En18
  input [18:0] Wgt_5_321, // sfix19_En18
  input [18:0] Wgt_5_322, // sfix19_En18
  input [18:0] Wgt_5_323, // sfix19_En18
  input [18:0] Wgt_5_324, // sfix19_En18
  input [18:0] Wgt_5_325, // sfix19_En18
  input [18:0] Wgt_5_326, // sfix19_En18
  input [18:0] Wgt_5_327, // sfix19_En18
  input [18:0] Wgt_5_328, // sfix19_En18
  input [18:0] Wgt_5_329, // sfix19_En18
  input [18:0] Wgt_5_330, // sfix19_En18
  input [18:0] Wgt_5_331, // sfix19_En18
  input [18:0] Wgt_5_332, // sfix19_En18
  input [18:0] Wgt_5_333, // sfix19_En18
  input [18:0] Wgt_5_334, // sfix19_En18
  input [18:0] Wgt_5_335, // sfix19_En18
  input [18:0] Wgt_5_336, // sfix19_En18
  input [18:0] Wgt_5_337, // sfix19_En18
  input [18:0] Wgt_5_338, // sfix19_En18
  input [18:0] Wgt_5_339, // sfix19_En18
  input [18:0] Wgt_5_340, // sfix19_En18
  input [18:0] Wgt_5_341, // sfix19_En18
  input [18:0] Wgt_5_342, // sfix19_En18
  input [18:0] Wgt_5_343, // sfix19_En18
  input [18:0] Wgt_5_344, // sfix19_En18
  input [18:0] Wgt_5_345, // sfix19_En18
  input [18:0] Wgt_5_346, // sfix19_En18
  input [18:0] Wgt_5_347, // sfix19_En18
  input [18:0] Wgt_5_348, // sfix19_En18
  input [18:0] Wgt_5_349, // sfix19_En18
  input [18:0] Wgt_5_350, // sfix19_En18
  input [18:0] Wgt_5_351, // sfix19_En18
  input [18:0] Wgt_5_352, // sfix19_En18
  input [18:0] Wgt_5_353, // sfix19_En18
  input [18:0] Wgt_5_354, // sfix19_En18
  input [18:0] Wgt_5_355, // sfix19_En18
  input [18:0] Wgt_5_356, // sfix19_En18
  input [18:0] Wgt_5_357, // sfix19_En18
  input [18:0] Wgt_5_358, // sfix19_En18
  input [18:0] Wgt_5_359, // sfix19_En18
  input [18:0] Wgt_5_360, // sfix19_En18
  input [18:0] Wgt_5_361, // sfix19_En18
  input [18:0] Wgt_5_362, // sfix19_En18
  input [18:0] Wgt_5_363, // sfix19_En18
  input [18:0] Wgt_5_364, // sfix19_En18
  input [18:0] Wgt_5_365, // sfix19_En18
  input [18:0] Wgt_5_366, // sfix19_En18
  input [18:0] Wgt_5_367, // sfix19_En18
  input [18:0] Wgt_5_368, // sfix19_En18
  input [18:0] Wgt_5_369, // sfix19_En18
  input [18:0] Wgt_5_370, // sfix19_En18
  input [18:0] Wgt_5_371, // sfix19_En18
  input [18:0] Wgt_5_372, // sfix19_En18
  input [18:0] Wgt_5_373, // sfix19_En18
  input [18:0] Wgt_5_374, // sfix19_En18
  input [18:0] Wgt_5_375, // sfix19_En18
  input [18:0] Wgt_5_376, // sfix19_En18
  input [18:0] Wgt_5_377, // sfix19_En18
  input [18:0] Wgt_5_378, // sfix19_En18
  input [18:0] Wgt_5_379, // sfix19_En18
  input [18:0] Wgt_5_380, // sfix19_En18
  input [18:0] Wgt_5_381, // sfix19_En18
  input [18:0] Wgt_5_382, // sfix19_En18
  input [18:0] Wgt_5_383, // sfix19_En18
  input [18:0] Wgt_5_384, // sfix19_En18
  input [18:0] Wgt_5_385, // sfix19_En18
  input [18:0] Wgt_5_386, // sfix19_En18
  input [18:0] Wgt_5_387, // sfix19_En18
  input [18:0] Wgt_5_388, // sfix19_En18
  input [18:0] Wgt_5_389, // sfix19_En18
  input [18:0] Wgt_5_390, // sfix19_En18
  input [18:0] Wgt_5_391, // sfix19_En18
  input [18:0] Wgt_5_392, // sfix19_En18
  input [18:0] Wgt_5_393, // sfix19_En18
  input [18:0] Wgt_5_394, // sfix19_En18
  input [18:0] Wgt_5_395, // sfix19_En18
  input [18:0] Wgt_5_396, // sfix19_En18
  input [18:0] Wgt_5_397, // sfix19_En18
  input [18:0] Wgt_5_398, // sfix19_En18
  input [18:0] Wgt_5_399, // sfix19_En18
  input [18:0] Wgt_5_400, // sfix19_En18
  input [18:0] Wgt_5_401, // sfix19_En18
  input [18:0] Wgt_5_402, // sfix19_En18
  input [18:0] Wgt_5_403, // sfix19_En18
  input [18:0] Wgt_5_404, // sfix19_En18
  input [18:0] Wgt_5_405, // sfix19_En18
  input [18:0] Wgt_5_406, // sfix19_En18
  input [18:0] Wgt_5_407, // sfix19_En18
  input [18:0] Wgt_5_408, // sfix19_En18
  input [18:0] Wgt_5_409, // sfix19_En18
  input [18:0] Wgt_5_410, // sfix19_En18
  input [18:0] Wgt_5_411, // sfix19_En18
  input [18:0] Wgt_5_412, // sfix19_En18
  input [18:0] Wgt_5_413, // sfix19_En18
  input [18:0] Wgt_5_414, // sfix19_En18
  input [18:0] Wgt_5_415, // sfix19_En18
  input [18:0] Wgt_5_416, // sfix19_En18
  input [18:0] Wgt_5_417, // sfix19_En18
  input [18:0] Wgt_5_418, // sfix19_En18
  input [18:0] Wgt_5_419, // sfix19_En18
  input [18:0] Wgt_5_420, // sfix19_En18
  input [18:0] Wgt_5_421, // sfix19_En18
  input [18:0] Wgt_5_422, // sfix19_En18
  input [18:0] Wgt_5_423, // sfix19_En18
  input [18:0] Wgt_5_424, // sfix19_En18
  input [18:0] Wgt_5_425, // sfix19_En18
  input [18:0] Wgt_5_426, // sfix19_En18
  input [18:0] Wgt_5_427, // sfix19_En18
  input [18:0] Wgt_5_428, // sfix19_En18
  input [18:0] Wgt_5_429, // sfix19_En18
  input [18:0] Wgt_5_430, // sfix19_En18
  input [18:0] Wgt_5_431, // sfix19_En18
  input [18:0] Wgt_5_432, // sfix19_En18
  input [18:0] Wgt_5_433, // sfix19_En18
  input [18:0] Wgt_5_434, // sfix19_En18
  input [18:0] Wgt_5_435, // sfix19_En18
  input [18:0] Wgt_5_436, // sfix19_En18
  input [18:0] Wgt_5_437, // sfix19_En18
  input [18:0] Wgt_5_438, // sfix19_En18
  input [18:0] Wgt_5_439, // sfix19_En18
  input [18:0] Wgt_5_440, // sfix19_En18
  input [18:0] Wgt_5_441, // sfix19_En18
  input [18:0] Wgt_5_442, // sfix19_En18
  input [18:0] Wgt_5_443, // sfix19_En18
  input [18:0] Wgt_5_444, // sfix19_En18
  input [18:0] Wgt_5_445, // sfix19_En18
  input [18:0] Wgt_5_446, // sfix19_En18
  input [18:0] Wgt_5_447, // sfix19_En18
  input [18:0] Wgt_5_448, // sfix19_En18
  input [18:0] Wgt_5_449, // sfix19_En18
  input [18:0] Wgt_5_450, // sfix19_En18
  input [18:0] Wgt_5_451, // sfix19_En18
  input [18:0] Wgt_5_452, // sfix19_En18
  input [18:0] Wgt_5_453, // sfix19_En18
  input [18:0] Wgt_5_454, // sfix19_En18
  input [18:0] Wgt_5_455, // sfix19_En18
  input [18:0] Wgt_5_456, // sfix19_En18
  input [18:0] Wgt_5_457, // sfix19_En18
  input [18:0] Wgt_5_458, // sfix19_En18
  input [18:0] Wgt_5_459, // sfix19_En18
  input [18:0] Wgt_5_460, // sfix19_En18
  input [18:0] Wgt_5_461, // sfix19_En18
  input [18:0] Wgt_5_462, // sfix19_En18
  input [18:0] Wgt_5_463, // sfix19_En18
  input [18:0] Wgt_5_464, // sfix19_En18
  input [18:0] Wgt_5_465, // sfix19_En18
  input [18:0] Wgt_5_466, // sfix19_En18
  input [18:0] Wgt_5_467, // sfix19_En18
  input [18:0] Wgt_5_468, // sfix19_En18
  input [18:0] Wgt_5_469, // sfix19_En18
  input [18:0] Wgt_5_470, // sfix19_En18
  input [18:0] Wgt_5_471, // sfix19_En18
  input [18:0] Wgt_5_472, // sfix19_En18
  input [18:0] Wgt_5_473, // sfix19_En18
  input [18:0] Wgt_5_474, // sfix19_En18
  input [18:0] Wgt_5_475, // sfix19_En18
  input [18:0] Wgt_5_476, // sfix19_En18
  input [18:0] Wgt_5_477, // sfix19_En18
  input [18:0] Wgt_5_478, // sfix19_En18
  input [18:0] Wgt_5_479, // sfix19_En18
  input [18:0] Wgt_5_480, // sfix19_En18
  input [18:0] Wgt_5_481, // sfix19_En18
  input [18:0] Wgt_5_482, // sfix19_En18
  input [18:0] Wgt_5_483, // sfix19_En18
  input [18:0] Wgt_5_484, // sfix19_En18
  input [18:0] Wgt_5_485, // sfix19_En18
  input [18:0] Wgt_5_486, // sfix19_En18
  input [18:0] Wgt_5_487, // sfix19_En18
  input [18:0] Wgt_5_488, // sfix19_En18
  input [18:0] Wgt_5_489, // sfix19_En18
  input [18:0] Wgt_5_490, // sfix19_En18
  input [18:0] Wgt_5_491, // sfix19_En18
  input [18:0] Wgt_5_492, // sfix19_En18
  input [18:0] Wgt_5_493, // sfix19_En18
  input [18:0] Wgt_5_494, // sfix19_En18
  input [18:0] Wgt_5_495, // sfix19_En18
  input [18:0] Wgt_5_496, // sfix19_En18
  input [18:0] Wgt_5_497, // sfix19_En18
  input [18:0] Wgt_5_498, // sfix19_En18
  input [18:0] Wgt_5_499, // sfix19_En18
  input [18:0] Wgt_5_500, // sfix19_En18
  input [18:0] Wgt_5_501, // sfix19_En18
  input [18:0] Wgt_5_502, // sfix19_En18
  input [18:0] Wgt_5_503, // sfix19_En18
  input [18:0] Wgt_5_504, // sfix19_En18
  input [18:0] Wgt_5_505, // sfix19_En18
  input [18:0] Wgt_5_506, // sfix19_En18
  input [18:0] Wgt_5_507, // sfix19_En18
  input [18:0] Wgt_5_508, // sfix19_En18
  input [18:0] Wgt_5_509, // sfix19_En18
  input [18:0] Wgt_5_510, // sfix19_En18
  input [18:0] Wgt_5_511, // sfix19_En18
  input [18:0] Wgt_5_512, // sfix19_En18
  input [18:0] Wgt_5_513, // sfix19_En18
  input [18:0] Wgt_5_514, // sfix19_En18
  input [18:0] Wgt_5_515, // sfix19_En18
  input [18:0] Wgt_5_516, // sfix19_En18
  input [18:0] Wgt_5_517, // sfix19_En18
  input [18:0] Wgt_5_518, // sfix19_En18
  input [18:0] Wgt_5_519, // sfix19_En18
  input [18:0] Wgt_5_520, // sfix19_En18
  input [18:0] Wgt_5_521, // sfix19_En18
  input [18:0] Wgt_5_522, // sfix19_En18
  input [18:0] Wgt_5_523, // sfix19_En18
  input [18:0] Wgt_5_524, // sfix19_En18
  input [18:0] Wgt_5_525, // sfix19_En18
  input [18:0] Wgt_5_526, // sfix19_En18
  input [18:0] Wgt_5_527, // sfix19_En18
  input [18:0] Wgt_5_528, // sfix19_En18
  input [18:0] Wgt_5_529, // sfix19_En18
  input [18:0] Wgt_5_530, // sfix19_En18
  input [18:0] Wgt_5_531, // sfix19_En18
  input [18:0] Wgt_5_532, // sfix19_En18
  input [18:0] Wgt_5_533, // sfix19_En18
  input [18:0] Wgt_5_534, // sfix19_En18
  input [18:0] Wgt_5_535, // sfix19_En18
  input [18:0] Wgt_5_536, // sfix19_En18
  input [18:0] Wgt_5_537, // sfix19_En18
  input [18:0] Wgt_5_538, // sfix19_En18
  input [18:0] Wgt_5_539, // sfix19_En18
  input [18:0] Wgt_5_540, // sfix19_En18
  input [18:0] Wgt_5_541, // sfix19_En18
  input [18:0] Wgt_5_542, // sfix19_En18
  input [18:0] Wgt_5_543, // sfix19_En18
  input [18:0] Wgt_5_544, // sfix19_En18
  input [18:0] Wgt_5_545, // sfix19_En18
  input [18:0] Wgt_5_546, // sfix19_En18
  input [18:0] Wgt_5_547, // sfix19_En18
  input [18:0] Wgt_5_548, // sfix19_En18
  input [18:0] Wgt_5_549, // sfix19_En18
  input [18:0] Wgt_5_550, // sfix19_En18
  input [18:0] Wgt_5_551, // sfix19_En18
  input [18:0] Wgt_5_552, // sfix19_En18
  input [18:0] Wgt_5_553, // sfix19_En18
  input [18:0] Wgt_5_554, // sfix19_En18
  input [18:0] Wgt_5_555, // sfix19_En18
  input [18:0] Wgt_5_556, // sfix19_En18
  input [18:0] Wgt_5_557, // sfix19_En18
  input [18:0] Wgt_5_558, // sfix19_En18
  input [18:0] Wgt_5_559, // sfix19_En18
  input [18:0] Wgt_5_560, // sfix19_En18
  input [18:0] Wgt_5_561, // sfix19_En18
  input [18:0] Wgt_5_562, // sfix19_En18
  input [18:0] Wgt_5_563, // sfix19_En18
  input [18:0] Wgt_5_564, // sfix19_En18
  input [18:0] Wgt_5_565, // sfix19_En18
  input [18:0] Wgt_5_566, // sfix19_En18
  input [18:0] Wgt_5_567, // sfix19_En18
  input [18:0] Wgt_5_568, // sfix19_En18
  input [18:0] Wgt_5_569, // sfix19_En18
  input [18:0] Wgt_5_570, // sfix19_En18
  input [18:0] Wgt_5_571, // sfix19_En18
  input [18:0] Wgt_5_572, // sfix19_En18
  input [18:0] Wgt_5_573, // sfix19_En18
  input [18:0] Wgt_5_574, // sfix19_En18
  input [18:0] Wgt_5_575, // sfix19_En18
  input [18:0] Wgt_5_576, // sfix19_En18
  input [18:0] Wgt_5_577, // sfix19_En18
  input [18:0] Wgt_5_578, // sfix19_En18
  input [18:0] Wgt_5_579, // sfix19_En18
  input [18:0] Wgt_5_580, // sfix19_En18
  input [18:0] Wgt_5_581, // sfix19_En18
  input [18:0] Wgt_5_582, // sfix19_En18
  input [18:0] Wgt_5_583, // sfix19_En18
  input [18:0] Wgt_5_584, // sfix19_En18
  input [18:0] Wgt_5_585, // sfix19_En18
  input [18:0] Wgt_5_586, // sfix19_En18
  input [18:0] Wgt_5_587, // sfix19_En18
  input [18:0] Wgt_5_588, // sfix19_En18
  input [18:0] Wgt_5_589, // sfix19_En18
  input [18:0] Wgt_5_590, // sfix19_En18
  input [18:0] Wgt_5_591, // sfix19_En18
  input [18:0] Wgt_5_592, // sfix19_En18
  input [18:0] Wgt_5_593, // sfix19_En18
  input [18:0] Wgt_5_594, // sfix19_En18
  input [18:0] Wgt_5_595, // sfix19_En18
  input [18:0] Wgt_5_596, // sfix19_En18
  input [18:0] Wgt_5_597, // sfix19_En18
  input [18:0] Wgt_5_598, // sfix19_En18
  input [18:0] Wgt_5_599, // sfix19_En18
  input [18:0] Wgt_5_600, // sfix19_En18
  input [18:0] Wgt_5_601, // sfix19_En18
  input [18:0] Wgt_5_602, // sfix19_En18
  input [18:0] Wgt_5_603, // sfix19_En18
  input [18:0] Wgt_5_604, // sfix19_En18
  input [18:0] Wgt_5_605, // sfix19_En18
  input [18:0] Wgt_5_606, // sfix19_En18
  input [18:0] Wgt_5_607, // sfix19_En18
  input [18:0] Wgt_5_608, // sfix19_En18
  input [18:0] Wgt_5_609, // sfix19_En18
  input [18:0] Wgt_5_610, // sfix19_En18
  input [18:0] Wgt_5_611, // sfix19_En18
  input [18:0] Wgt_5_612, // sfix19_En18
  input [18:0] Wgt_5_613, // sfix19_En18
  input [18:0] Wgt_5_614, // sfix19_En18
  input [18:0] Wgt_5_615, // sfix19_En18
  input [18:0] Wgt_5_616, // sfix19_En18
  input [18:0] Wgt_5_617, // sfix19_En18
  input [18:0] Wgt_5_618, // sfix19_En18
  input [18:0] Wgt_5_619, // sfix19_En18
  input [18:0] Wgt_5_620, // sfix19_En18
  input [18:0] Wgt_5_621, // sfix19_En18
  input [18:0] Wgt_5_622, // sfix19_En18
  input [18:0] Wgt_5_623, // sfix19_En18
  input [18:0] Wgt_5_624, // sfix19_En18
  input [18:0] Wgt_5_625, // sfix19_En18
  input [18:0] Wgt_5_626, // sfix19_En18
  input [18:0] Wgt_5_627, // sfix19_En18
  input [18:0] Wgt_5_628, // sfix19_En18
  input [18:0] Wgt_5_629, // sfix19_En18
  input [18:0] Wgt_5_630, // sfix19_En18
  input [18:0] Wgt_5_631, // sfix19_En18
  input [18:0] Wgt_5_632, // sfix19_En18
  input [18:0] Wgt_5_633, // sfix19_En18
  input [18:0] Wgt_5_634, // sfix19_En18
  input [18:0] Wgt_5_635, // sfix19_En18
  input [18:0] Wgt_5_636, // sfix19_En18
  input [18:0] Wgt_5_637, // sfix19_En18
  input [18:0] Wgt_5_638, // sfix19_En18
  input [18:0] Wgt_5_639, // sfix19_En18
  input [18:0] Wgt_5_640, // sfix19_En18
  input [18:0] Wgt_5_641, // sfix19_En18
  input [18:0] Wgt_5_642, // sfix19_En18
  input [18:0] Wgt_5_643, // sfix19_En18
  input [18:0] Wgt_5_644, // sfix19_En18
  input [18:0] Wgt_5_645, // sfix19_En18
  input [18:0] Wgt_5_646, // sfix19_En18
  input [18:0] Wgt_5_647, // sfix19_En18
  input [18:0] Wgt_5_648, // sfix19_En18
  input [18:0] Wgt_5_649, // sfix19_En18
  input [18:0] Wgt_5_650, // sfix19_En18
  input [18:0] Wgt_5_651, // sfix19_En18
  input [18:0] Wgt_5_652, // sfix19_En18
  input [18:0] Wgt_5_653, // sfix19_En18
  input [18:0] Wgt_5_654, // sfix19_En18
  input [18:0] Wgt_5_655, // sfix19_En18
  input [18:0] Wgt_5_656, // sfix19_En18
  input [18:0] Wgt_5_657, // sfix19_En18
  input [18:0] Wgt_5_658, // sfix19_En18
  input [18:0] Wgt_5_659, // sfix19_En18
  input [18:0] Wgt_5_660, // sfix19_En18
  input [18:0] Wgt_5_661, // sfix19_En18
  input [18:0] Wgt_5_662, // sfix19_En18
  input [18:0] Wgt_5_663, // sfix19_En18
  input [18:0] Wgt_5_664, // sfix19_En18
  input [18:0] Wgt_5_665, // sfix19_En18
  input [18:0] Wgt_5_666, // sfix19_En18
  input [18:0] Wgt_5_667, // sfix19_En18
  input [18:0] Wgt_5_668, // sfix19_En18
  input [18:0] Wgt_5_669, // sfix19_En18
  input [18:0] Wgt_5_670, // sfix19_En18
  input [18:0] Wgt_5_671, // sfix19_En18
  input [18:0] Wgt_5_672, // sfix19_En18
  input [18:0] Wgt_5_673, // sfix19_En18
  input [18:0] Wgt_5_674, // sfix19_En18
  input [18:0] Wgt_5_675, // sfix19_En18
  input [18:0] Wgt_5_676, // sfix19_En18
  input [18:0] Wgt_5_677, // sfix19_En18
  input [18:0] Wgt_5_678, // sfix19_En18
  input [18:0] Wgt_5_679, // sfix19_En18
  input [18:0] Wgt_5_680, // sfix19_En18
  input [18:0] Wgt_5_681, // sfix19_En18
  input [18:0] Wgt_5_682, // sfix19_En18
  input [18:0] Wgt_5_683, // sfix19_En18
  input [18:0] Wgt_5_684, // sfix19_En18
  input [18:0] Wgt_5_685, // sfix19_En18
  input [18:0] Wgt_5_686, // sfix19_En18
  input [18:0] Wgt_5_687, // sfix19_En18
  input [18:0] Wgt_5_688, // sfix19_En18
  input [18:0] Wgt_5_689, // sfix19_En18
  input [18:0] Wgt_5_690, // sfix19_En18
  input [18:0] Wgt_5_691, // sfix19_En18
  input [18:0] Wgt_5_692, // sfix19_En18
  input [18:0] Wgt_5_693, // sfix19_En18
  input [18:0] Wgt_5_694, // sfix19_En18
  input [18:0] Wgt_5_695, // sfix19_En18
  input [18:0] Wgt_5_696, // sfix19_En18
  input [18:0] Wgt_5_697, // sfix19_En18
  input [18:0] Wgt_5_698, // sfix19_En18
  input [18:0] Wgt_5_699, // sfix19_En18
  input [18:0] Wgt_5_700, // sfix19_En18
  input [18:0] Wgt_5_701, // sfix19_En18
  input [18:0] Wgt_5_702, // sfix19_En18
  input [18:0] Wgt_5_703, // sfix19_En18
  input [18:0] Wgt_5_704, // sfix19_En18
  input [18:0] Wgt_5_705, // sfix19_En18
  input [18:0] Wgt_5_706, // sfix19_En18
  input [18:0] Wgt_5_707, // sfix19_En18
  input [18:0] Wgt_5_708, // sfix19_En18
  input [18:0] Wgt_5_709, // sfix19_En18
  input [18:0] Wgt_5_710, // sfix19_En18
  input [18:0] Wgt_5_711, // sfix19_En18
  input [18:0] Wgt_5_712, // sfix19_En18
  input [18:0] Wgt_5_713, // sfix19_En18
  input [18:0] Wgt_5_714, // sfix19_En18
  input [18:0] Wgt_5_715, // sfix19_En18
  input [18:0] Wgt_5_716, // sfix19_En18
  input [18:0] Wgt_5_717, // sfix19_En18
  input [18:0] Wgt_5_718, // sfix19_En18
  input [18:0] Wgt_5_719, // sfix19_En18
  input [18:0] Wgt_5_720, // sfix19_En18
  input [18:0] Wgt_5_721, // sfix19_En18
  input [18:0] Wgt_5_722, // sfix19_En18
  input [18:0] Wgt_5_723, // sfix19_En18
  input [18:0] Wgt_5_724, // sfix19_En18
  input [18:0] Wgt_5_725, // sfix19_En18
  input [18:0] Wgt_5_726, // sfix19_En18
  input [18:0] Wgt_5_727, // sfix19_En18
  input [18:0] Wgt_5_728, // sfix19_En18
  input [18:0] Wgt_5_729, // sfix19_En18
  input [18:0] Wgt_5_730, // sfix19_En18
  input [18:0] Wgt_5_731, // sfix19_En18
  input [18:0] Wgt_5_732, // sfix19_En18
  input [18:0] Wgt_5_733, // sfix19_En18
  input [18:0] Wgt_5_734, // sfix19_En18
  input [18:0] Wgt_5_735, // sfix19_En18
  input [18:0] Wgt_5_736, // sfix19_En18
  input [18:0] Wgt_5_737, // sfix19_En18
  input [18:0] Wgt_5_738, // sfix19_En18
  input [18:0] Wgt_5_739, // sfix19_En18
  input [18:0] Wgt_5_740, // sfix19_En18
  input [18:0] Wgt_5_741, // sfix19_En18
  input [18:0] Wgt_5_742, // sfix19_En18
  input [18:0] Wgt_5_743, // sfix19_En18
  input [18:0] Wgt_5_744, // sfix19_En18
  input [18:0] Wgt_5_745, // sfix19_En18
  input [18:0] Wgt_5_746, // sfix19_En18
  input [18:0] Wgt_5_747, // sfix19_En18
  input [18:0] Wgt_5_748, // sfix19_En18
  input [18:0] Wgt_5_749, // sfix19_En18
  input [18:0] Wgt_5_750, // sfix19_En18
  input [18:0] Wgt_5_751, // sfix19_En18
  input [18:0] Wgt_5_752, // sfix19_En18
  input [18:0] Wgt_5_753, // sfix19_En18
  input [18:0] Wgt_5_754, // sfix19_En18
  input [18:0] Wgt_5_755, // sfix19_En18
  input [18:0] Wgt_5_756, // sfix19_En18
  input [18:0] Wgt_5_757, // sfix19_En18
  input [18:0] Wgt_5_758, // sfix19_En18
  input [18:0] Wgt_5_759, // sfix19_En18
  input [18:0] Wgt_5_760, // sfix19_En18
  input [18:0] Wgt_5_761, // sfix19_En18
  input [18:0] Wgt_5_762, // sfix19_En18
  input [18:0] Wgt_5_763, // sfix19_En18
  input [18:0] Wgt_5_764, // sfix19_En18
  input [18:0] Wgt_5_765, // sfix19_En18
  input [18:0] Wgt_5_766, // sfix19_En18
  input [18:0] Wgt_5_767, // sfix19_En18
  input [18:0] Wgt_5_768, // sfix19_En18
  input [18:0] Wgt_5_769, // sfix19_En18
  input [18:0] Wgt_5_770, // sfix19_En18
  input [18:0] Wgt_5_771, // sfix19_En18
  input [18:0] Wgt_5_772, // sfix19_En18
  input [18:0] Wgt_5_773, // sfix19_En18
  input [18:0] Wgt_5_774, // sfix19_En18
  input [18:0] Wgt_5_775, // sfix19_En18
  input [18:0] Wgt_5_776, // sfix19_En18
  input [18:0] Wgt_5_777, // sfix19_En18
  input [18:0] Wgt_5_778, // sfix19_En18
  input [18:0] Wgt_5_779, // sfix19_En18
  input [18:0] Wgt_5_780, // sfix19_En18
  input [18:0] Wgt_5_781, // sfix19_En18
  input [18:0] Wgt_5_782, // sfix19_En18
  input [18:0] Wgt_5_783, // sfix19_En18
  input [18:0] Wgt_5_784, // sfix19_En18
  input [18:0] Wgt_6_0, // sfix19_En18
  input [18:0] Wgt_6_1, // sfix19_En18
  input [18:0] Wgt_6_2, // sfix19_En18
  input [18:0] Wgt_6_3, // sfix19_En18
  input [18:0] Wgt_6_4, // sfix19_En18
  input [18:0] Wgt_6_5, // sfix19_En18
  input [18:0] Wgt_6_6, // sfix19_En18
  input [18:0] Wgt_6_7, // sfix19_En18
  input [18:0] Wgt_6_8, // sfix19_En18
  input [18:0] Wgt_6_9, // sfix19_En18
  input [18:0] Wgt_6_10, // sfix19_En18
  input [18:0] Wgt_6_11, // sfix19_En18
  input [18:0] Wgt_6_12, // sfix19_En18
  input [18:0] Wgt_6_13, // sfix19_En18
  input [18:0] Wgt_6_14, // sfix19_En18
  input [18:0] Wgt_6_15, // sfix19_En18
  input [18:0] Wgt_6_16, // sfix19_En18
  input [18:0] Wgt_6_17, // sfix19_En18
  input [18:0] Wgt_6_18, // sfix19_En18
  input [18:0] Wgt_6_19, // sfix19_En18
  input [18:0] Wgt_6_20, // sfix19_En18
  input [18:0] Wgt_6_21, // sfix19_En18
  input [18:0] Wgt_6_22, // sfix19_En18
  input [18:0] Wgt_6_23, // sfix19_En18
  input [18:0] Wgt_6_24, // sfix19_En18
  input [18:0] Wgt_6_25, // sfix19_En18
  input [18:0] Wgt_6_26, // sfix19_En18
  input [18:0] Wgt_6_27, // sfix19_En18
  input [18:0] Wgt_6_28, // sfix19_En18
  input [18:0] Wgt_6_29, // sfix19_En18
  input [18:0] Wgt_6_30, // sfix19_En18
  input [18:0] Wgt_6_31, // sfix19_En18
  input [18:0] Wgt_6_32, // sfix19_En18
  input [18:0] Wgt_6_33, // sfix19_En18
  input [18:0] Wgt_6_34, // sfix19_En18
  input [18:0] Wgt_6_35, // sfix19_En18
  input [18:0] Wgt_6_36, // sfix19_En18
  input [18:0] Wgt_6_37, // sfix19_En18
  input [18:0] Wgt_6_38, // sfix19_En18
  input [18:0] Wgt_6_39, // sfix19_En18
  input [18:0] Wgt_6_40, // sfix19_En18
  input [18:0] Wgt_6_41, // sfix19_En18
  input [18:0] Wgt_6_42, // sfix19_En18
  input [18:0] Wgt_6_43, // sfix19_En18
  input [18:0] Wgt_6_44, // sfix19_En18
  input [18:0] Wgt_6_45, // sfix19_En18
  input [18:0] Wgt_6_46, // sfix19_En18
  input [18:0] Wgt_6_47, // sfix19_En18
  input [18:0] Wgt_6_48, // sfix19_En18
  input [18:0] Wgt_6_49, // sfix19_En18
  input [18:0] Wgt_6_50, // sfix19_En18
  input [18:0] Wgt_6_51, // sfix19_En18
  input [18:0] Wgt_6_52, // sfix19_En18
  input [18:0] Wgt_6_53, // sfix19_En18
  input [18:0] Wgt_6_54, // sfix19_En18
  input [18:0] Wgt_6_55, // sfix19_En18
  input [18:0] Wgt_6_56, // sfix19_En18
  input [18:0] Wgt_6_57, // sfix19_En18
  input [18:0] Wgt_6_58, // sfix19_En18
  input [18:0] Wgt_6_59, // sfix19_En18
  input [18:0] Wgt_6_60, // sfix19_En18
  input [18:0] Wgt_6_61, // sfix19_En18
  input [18:0] Wgt_6_62, // sfix19_En18
  input [18:0] Wgt_6_63, // sfix19_En18
  input [18:0] Wgt_6_64, // sfix19_En18
  input [18:0] Wgt_6_65, // sfix19_En18
  input [18:0] Wgt_6_66, // sfix19_En18
  input [18:0] Wgt_6_67, // sfix19_En18
  input [18:0] Wgt_6_68, // sfix19_En18
  input [18:0] Wgt_6_69, // sfix19_En18
  input [18:0] Wgt_6_70, // sfix19_En18
  input [18:0] Wgt_6_71, // sfix19_En18
  input [18:0] Wgt_6_72, // sfix19_En18
  input [18:0] Wgt_6_73, // sfix19_En18
  input [18:0] Wgt_6_74, // sfix19_En18
  input [18:0] Wgt_6_75, // sfix19_En18
  input [18:0] Wgt_6_76, // sfix19_En18
  input [18:0] Wgt_6_77, // sfix19_En18
  input [18:0] Wgt_6_78, // sfix19_En18
  input [18:0] Wgt_6_79, // sfix19_En18
  input [18:0] Wgt_6_80, // sfix19_En18
  input [18:0] Wgt_6_81, // sfix19_En18
  input [18:0] Wgt_6_82, // sfix19_En18
  input [18:0] Wgt_6_83, // sfix19_En18
  input [18:0] Wgt_6_84, // sfix19_En18
  input [18:0] Wgt_6_85, // sfix19_En18
  input [18:0] Wgt_6_86, // sfix19_En18
  input [18:0] Wgt_6_87, // sfix19_En18
  input [18:0] Wgt_6_88, // sfix19_En18
  input [18:0] Wgt_6_89, // sfix19_En18
  input [18:0] Wgt_6_90, // sfix19_En18
  input [18:0] Wgt_6_91, // sfix19_En18
  input [18:0] Wgt_6_92, // sfix19_En18
  input [18:0] Wgt_6_93, // sfix19_En18
  input [18:0] Wgt_6_94, // sfix19_En18
  input [18:0] Wgt_6_95, // sfix19_En18
  input [18:0] Wgt_6_96, // sfix19_En18
  input [18:0] Wgt_6_97, // sfix19_En18
  input [18:0] Wgt_6_98, // sfix19_En18
  input [18:0] Wgt_6_99, // sfix19_En18
  input [18:0] Wgt_6_100, // sfix19_En18
  input [18:0] Wgt_6_101, // sfix19_En18
  input [18:0] Wgt_6_102, // sfix19_En18
  input [18:0] Wgt_6_103, // sfix19_En18
  input [18:0] Wgt_6_104, // sfix19_En18
  input [18:0] Wgt_6_105, // sfix19_En18
  input [18:0] Wgt_6_106, // sfix19_En18
  input [18:0] Wgt_6_107, // sfix19_En18
  input [18:0] Wgt_6_108, // sfix19_En18
  input [18:0] Wgt_6_109, // sfix19_En18
  input [18:0] Wgt_6_110, // sfix19_En18
  input [18:0] Wgt_6_111, // sfix19_En18
  input [18:0] Wgt_6_112, // sfix19_En18
  input [18:0] Wgt_6_113, // sfix19_En18
  input [18:0] Wgt_6_114, // sfix19_En18
  input [18:0] Wgt_6_115, // sfix19_En18
  input [18:0] Wgt_6_116, // sfix19_En18
  input [18:0] Wgt_6_117, // sfix19_En18
  input [18:0] Wgt_6_118, // sfix19_En18
  input [18:0] Wgt_6_119, // sfix19_En18
  input [18:0] Wgt_6_120, // sfix19_En18
  input [18:0] Wgt_6_121, // sfix19_En18
  input [18:0] Wgt_6_122, // sfix19_En18
  input [18:0] Wgt_6_123, // sfix19_En18
  input [18:0] Wgt_6_124, // sfix19_En18
  input [18:0] Wgt_6_125, // sfix19_En18
  input [18:0] Wgt_6_126, // sfix19_En18
  input [18:0] Wgt_6_127, // sfix19_En18
  input [18:0] Wgt_6_128, // sfix19_En18
  input [18:0] Wgt_6_129, // sfix19_En18
  input [18:0] Wgt_6_130, // sfix19_En18
  input [18:0] Wgt_6_131, // sfix19_En18
  input [18:0] Wgt_6_132, // sfix19_En18
  input [18:0] Wgt_6_133, // sfix19_En18
  input [18:0] Wgt_6_134, // sfix19_En18
  input [18:0] Wgt_6_135, // sfix19_En18
  input [18:0] Wgt_6_136, // sfix19_En18
  input [18:0] Wgt_6_137, // sfix19_En18
  input [18:0] Wgt_6_138, // sfix19_En18
  input [18:0] Wgt_6_139, // sfix19_En18
  input [18:0] Wgt_6_140, // sfix19_En18
  input [18:0] Wgt_6_141, // sfix19_En18
  input [18:0] Wgt_6_142, // sfix19_En18
  input [18:0] Wgt_6_143, // sfix19_En18
  input [18:0] Wgt_6_144, // sfix19_En18
  input [18:0] Wgt_6_145, // sfix19_En18
  input [18:0] Wgt_6_146, // sfix19_En18
  input [18:0] Wgt_6_147, // sfix19_En18
  input [18:0] Wgt_6_148, // sfix19_En18
  input [18:0] Wgt_6_149, // sfix19_En18
  input [18:0] Wgt_6_150, // sfix19_En18
  input [18:0] Wgt_6_151, // sfix19_En18
  input [18:0] Wgt_6_152, // sfix19_En18
  input [18:0] Wgt_6_153, // sfix19_En18
  input [18:0] Wgt_6_154, // sfix19_En18
  input [18:0] Wgt_6_155, // sfix19_En18
  input [18:0] Wgt_6_156, // sfix19_En18
  input [18:0] Wgt_6_157, // sfix19_En18
  input [18:0] Wgt_6_158, // sfix19_En18
  input [18:0] Wgt_6_159, // sfix19_En18
  input [18:0] Wgt_6_160, // sfix19_En18
  input [18:0] Wgt_6_161, // sfix19_En18
  input [18:0] Wgt_6_162, // sfix19_En18
  input [18:0] Wgt_6_163, // sfix19_En18
  input [18:0] Wgt_6_164, // sfix19_En18
  input [18:0] Wgt_6_165, // sfix19_En18
  input [18:0] Wgt_6_166, // sfix19_En18
  input [18:0] Wgt_6_167, // sfix19_En18
  input [18:0] Wgt_6_168, // sfix19_En18
  input [18:0] Wgt_6_169, // sfix19_En18
  input [18:0] Wgt_6_170, // sfix19_En18
  input [18:0] Wgt_6_171, // sfix19_En18
  input [18:0] Wgt_6_172, // sfix19_En18
  input [18:0] Wgt_6_173, // sfix19_En18
  input [18:0] Wgt_6_174, // sfix19_En18
  input [18:0] Wgt_6_175, // sfix19_En18
  input [18:0] Wgt_6_176, // sfix19_En18
  input [18:0] Wgt_6_177, // sfix19_En18
  input [18:0] Wgt_6_178, // sfix19_En18
  input [18:0] Wgt_6_179, // sfix19_En18
  input [18:0] Wgt_6_180, // sfix19_En18
  input [18:0] Wgt_6_181, // sfix19_En18
  input [18:0] Wgt_6_182, // sfix19_En18
  input [18:0] Wgt_6_183, // sfix19_En18
  input [18:0] Wgt_6_184, // sfix19_En18
  input [18:0] Wgt_6_185, // sfix19_En18
  input [18:0] Wgt_6_186, // sfix19_En18
  input [18:0] Wgt_6_187, // sfix19_En18
  input [18:0] Wgt_6_188, // sfix19_En18
  input [18:0] Wgt_6_189, // sfix19_En18
  input [18:0] Wgt_6_190, // sfix19_En18
  input [18:0] Wgt_6_191, // sfix19_En18
  input [18:0] Wgt_6_192, // sfix19_En18
  input [18:0] Wgt_6_193, // sfix19_En18
  input [18:0] Wgt_6_194, // sfix19_En18
  input [18:0] Wgt_6_195, // sfix19_En18
  input [18:0] Wgt_6_196, // sfix19_En18
  input [18:0] Wgt_6_197, // sfix19_En18
  input [18:0] Wgt_6_198, // sfix19_En18
  input [18:0] Wgt_6_199, // sfix19_En18
  input [18:0] Wgt_6_200, // sfix19_En18
  input [18:0] Wgt_6_201, // sfix19_En18
  input [18:0] Wgt_6_202, // sfix19_En18
  input [18:0] Wgt_6_203, // sfix19_En18
  input [18:0] Wgt_6_204, // sfix19_En18
  input [18:0] Wgt_6_205, // sfix19_En18
  input [18:0] Wgt_6_206, // sfix19_En18
  input [18:0] Wgt_6_207, // sfix19_En18
  input [18:0] Wgt_6_208, // sfix19_En18
  input [18:0] Wgt_6_209, // sfix19_En18
  input [18:0] Wgt_6_210, // sfix19_En18
  input [18:0] Wgt_6_211, // sfix19_En18
  input [18:0] Wgt_6_212, // sfix19_En18
  input [18:0] Wgt_6_213, // sfix19_En18
  input [18:0] Wgt_6_214, // sfix19_En18
  input [18:0] Wgt_6_215, // sfix19_En18
  input [18:0] Wgt_6_216, // sfix19_En18
  input [18:0] Wgt_6_217, // sfix19_En18
  input [18:0] Wgt_6_218, // sfix19_En18
  input [18:0] Wgt_6_219, // sfix19_En18
  input [18:0] Wgt_6_220, // sfix19_En18
  input [18:0] Wgt_6_221, // sfix19_En18
  input [18:0] Wgt_6_222, // sfix19_En18
  input [18:0] Wgt_6_223, // sfix19_En18
  input [18:0] Wgt_6_224, // sfix19_En18
  input [18:0] Wgt_6_225, // sfix19_En18
  input [18:0] Wgt_6_226, // sfix19_En18
  input [18:0] Wgt_6_227, // sfix19_En18
  input [18:0] Wgt_6_228, // sfix19_En18
  input [18:0] Wgt_6_229, // sfix19_En18
  input [18:0] Wgt_6_230, // sfix19_En18
  input [18:0] Wgt_6_231, // sfix19_En18
  input [18:0] Wgt_6_232, // sfix19_En18
  input [18:0] Wgt_6_233, // sfix19_En18
  input [18:0] Wgt_6_234, // sfix19_En18
  input [18:0] Wgt_6_235, // sfix19_En18
  input [18:0] Wgt_6_236, // sfix19_En18
  input [18:0] Wgt_6_237, // sfix19_En18
  input [18:0] Wgt_6_238, // sfix19_En18
  input [18:0] Wgt_6_239, // sfix19_En18
  input [18:0] Wgt_6_240, // sfix19_En18
  input [18:0] Wgt_6_241, // sfix19_En18
  input [18:0] Wgt_6_242, // sfix19_En18
  input [18:0] Wgt_6_243, // sfix19_En18
  input [18:0] Wgt_6_244, // sfix19_En18
  input [18:0] Wgt_6_245, // sfix19_En18
  input [18:0] Wgt_6_246, // sfix19_En18
  input [18:0] Wgt_6_247, // sfix19_En18
  input [18:0] Wgt_6_248, // sfix19_En18
  input [18:0] Wgt_6_249, // sfix19_En18
  input [18:0] Wgt_6_250, // sfix19_En18
  input [18:0] Wgt_6_251, // sfix19_En18
  input [18:0] Wgt_6_252, // sfix19_En18
  input [18:0] Wgt_6_253, // sfix19_En18
  input [18:0] Wgt_6_254, // sfix19_En18
  input [18:0] Wgt_6_255, // sfix19_En18
  input [18:0] Wgt_6_256, // sfix19_En18
  input [18:0] Wgt_6_257, // sfix19_En18
  input [18:0] Wgt_6_258, // sfix19_En18
  input [18:0] Wgt_6_259, // sfix19_En18
  input [18:0] Wgt_6_260, // sfix19_En18
  input [18:0] Wgt_6_261, // sfix19_En18
  input [18:0] Wgt_6_262, // sfix19_En18
  input [18:0] Wgt_6_263, // sfix19_En18
  input [18:0] Wgt_6_264, // sfix19_En18
  input [18:0] Wgt_6_265, // sfix19_En18
  input [18:0] Wgt_6_266, // sfix19_En18
  input [18:0] Wgt_6_267, // sfix19_En18
  input [18:0] Wgt_6_268, // sfix19_En18
  input [18:0] Wgt_6_269, // sfix19_En18
  input [18:0] Wgt_6_270, // sfix19_En18
  input [18:0] Wgt_6_271, // sfix19_En18
  input [18:0] Wgt_6_272, // sfix19_En18
  input [18:0] Wgt_6_273, // sfix19_En18
  input [18:0] Wgt_6_274, // sfix19_En18
  input [18:0] Wgt_6_275, // sfix19_En18
  input [18:0] Wgt_6_276, // sfix19_En18
  input [18:0] Wgt_6_277, // sfix19_En18
  input [18:0] Wgt_6_278, // sfix19_En18
  input [18:0] Wgt_6_279, // sfix19_En18
  input [18:0] Wgt_6_280, // sfix19_En18
  input [18:0] Wgt_6_281, // sfix19_En18
  input [18:0] Wgt_6_282, // sfix19_En18
  input [18:0] Wgt_6_283, // sfix19_En18
  input [18:0] Wgt_6_284, // sfix19_En18
  input [18:0] Wgt_6_285, // sfix19_En18
  input [18:0] Wgt_6_286, // sfix19_En18
  input [18:0] Wgt_6_287, // sfix19_En18
  input [18:0] Wgt_6_288, // sfix19_En18
  input [18:0] Wgt_6_289, // sfix19_En18
  input [18:0] Wgt_6_290, // sfix19_En18
  input [18:0] Wgt_6_291, // sfix19_En18
  input [18:0] Wgt_6_292, // sfix19_En18
  input [18:0] Wgt_6_293, // sfix19_En18
  input [18:0] Wgt_6_294, // sfix19_En18
  input [18:0] Wgt_6_295, // sfix19_En18
  input [18:0] Wgt_6_296, // sfix19_En18
  input [18:0] Wgt_6_297, // sfix19_En18
  input [18:0] Wgt_6_298, // sfix19_En18
  input [18:0] Wgt_6_299, // sfix19_En18
  input [18:0] Wgt_6_300, // sfix19_En18
  input [18:0] Wgt_6_301, // sfix19_En18
  input [18:0] Wgt_6_302, // sfix19_En18
  input [18:0] Wgt_6_303, // sfix19_En18
  input [18:0] Wgt_6_304, // sfix19_En18
  input [18:0] Wgt_6_305, // sfix19_En18
  input [18:0] Wgt_6_306, // sfix19_En18
  input [18:0] Wgt_6_307, // sfix19_En18
  input [18:0] Wgt_6_308, // sfix19_En18
  input [18:0] Wgt_6_309, // sfix19_En18
  input [18:0] Wgt_6_310, // sfix19_En18
  input [18:0] Wgt_6_311, // sfix19_En18
  input [18:0] Wgt_6_312, // sfix19_En18
  input [18:0] Wgt_6_313, // sfix19_En18
  input [18:0] Wgt_6_314, // sfix19_En18
  input [18:0] Wgt_6_315, // sfix19_En18
  input [18:0] Wgt_6_316, // sfix19_En18
  input [18:0] Wgt_6_317, // sfix19_En18
  input [18:0] Wgt_6_318, // sfix19_En18
  input [18:0] Wgt_6_319, // sfix19_En18
  input [18:0] Wgt_6_320, // sfix19_En18
  input [18:0] Wgt_6_321, // sfix19_En18
  input [18:0] Wgt_6_322, // sfix19_En18
  input [18:0] Wgt_6_323, // sfix19_En18
  input [18:0] Wgt_6_324, // sfix19_En18
  input [18:0] Wgt_6_325, // sfix19_En18
  input [18:0] Wgt_6_326, // sfix19_En18
  input [18:0] Wgt_6_327, // sfix19_En18
  input [18:0] Wgt_6_328, // sfix19_En18
  input [18:0] Wgt_6_329, // sfix19_En18
  input [18:0] Wgt_6_330, // sfix19_En18
  input [18:0] Wgt_6_331, // sfix19_En18
  input [18:0] Wgt_6_332, // sfix19_En18
  input [18:0] Wgt_6_333, // sfix19_En18
  input [18:0] Wgt_6_334, // sfix19_En18
  input [18:0] Wgt_6_335, // sfix19_En18
  input [18:0] Wgt_6_336, // sfix19_En18
  input [18:0] Wgt_6_337, // sfix19_En18
  input [18:0] Wgt_6_338, // sfix19_En18
  input [18:0] Wgt_6_339, // sfix19_En18
  input [18:0] Wgt_6_340, // sfix19_En18
  input [18:0] Wgt_6_341, // sfix19_En18
  input [18:0] Wgt_6_342, // sfix19_En18
  input [18:0] Wgt_6_343, // sfix19_En18
  input [18:0] Wgt_6_344, // sfix19_En18
  input [18:0] Wgt_6_345, // sfix19_En18
  input [18:0] Wgt_6_346, // sfix19_En18
  input [18:0] Wgt_6_347, // sfix19_En18
  input [18:0] Wgt_6_348, // sfix19_En18
  input [18:0] Wgt_6_349, // sfix19_En18
  input [18:0] Wgt_6_350, // sfix19_En18
  input [18:0] Wgt_6_351, // sfix19_En18
  input [18:0] Wgt_6_352, // sfix19_En18
  input [18:0] Wgt_6_353, // sfix19_En18
  input [18:0] Wgt_6_354, // sfix19_En18
  input [18:0] Wgt_6_355, // sfix19_En18
  input [18:0] Wgt_6_356, // sfix19_En18
  input [18:0] Wgt_6_357, // sfix19_En18
  input [18:0] Wgt_6_358, // sfix19_En18
  input [18:0] Wgt_6_359, // sfix19_En18
  input [18:0] Wgt_6_360, // sfix19_En18
  input [18:0] Wgt_6_361, // sfix19_En18
  input [18:0] Wgt_6_362, // sfix19_En18
  input [18:0] Wgt_6_363, // sfix19_En18
  input [18:0] Wgt_6_364, // sfix19_En18
  input [18:0] Wgt_6_365, // sfix19_En18
  input [18:0] Wgt_6_366, // sfix19_En18
  input [18:0] Wgt_6_367, // sfix19_En18
  input [18:0] Wgt_6_368, // sfix19_En18
  input [18:0] Wgt_6_369, // sfix19_En18
  input [18:0] Wgt_6_370, // sfix19_En18
  input [18:0] Wgt_6_371, // sfix19_En18
  input [18:0] Wgt_6_372, // sfix19_En18
  input [18:0] Wgt_6_373, // sfix19_En18
  input [18:0] Wgt_6_374, // sfix19_En18
  input [18:0] Wgt_6_375, // sfix19_En18
  input [18:0] Wgt_6_376, // sfix19_En18
  input [18:0] Wgt_6_377, // sfix19_En18
  input [18:0] Wgt_6_378, // sfix19_En18
  input [18:0] Wgt_6_379, // sfix19_En18
  input [18:0] Wgt_6_380, // sfix19_En18
  input [18:0] Wgt_6_381, // sfix19_En18
  input [18:0] Wgt_6_382, // sfix19_En18
  input [18:0] Wgt_6_383, // sfix19_En18
  input [18:0] Wgt_6_384, // sfix19_En18
  input [18:0] Wgt_6_385, // sfix19_En18
  input [18:0] Wgt_6_386, // sfix19_En18
  input [18:0] Wgt_6_387, // sfix19_En18
  input [18:0] Wgt_6_388, // sfix19_En18
  input [18:0] Wgt_6_389, // sfix19_En18
  input [18:0] Wgt_6_390, // sfix19_En18
  input [18:0] Wgt_6_391, // sfix19_En18
  input [18:0] Wgt_6_392, // sfix19_En18
  input [18:0] Wgt_6_393, // sfix19_En18
  input [18:0] Wgt_6_394, // sfix19_En18
  input [18:0] Wgt_6_395, // sfix19_En18
  input [18:0] Wgt_6_396, // sfix19_En18
  input [18:0] Wgt_6_397, // sfix19_En18
  input [18:0] Wgt_6_398, // sfix19_En18
  input [18:0] Wgt_6_399, // sfix19_En18
  input [18:0] Wgt_6_400, // sfix19_En18
  input [18:0] Wgt_6_401, // sfix19_En18
  input [18:0] Wgt_6_402, // sfix19_En18
  input [18:0] Wgt_6_403, // sfix19_En18
  input [18:0] Wgt_6_404, // sfix19_En18
  input [18:0] Wgt_6_405, // sfix19_En18
  input [18:0] Wgt_6_406, // sfix19_En18
  input [18:0] Wgt_6_407, // sfix19_En18
  input [18:0] Wgt_6_408, // sfix19_En18
  input [18:0] Wgt_6_409, // sfix19_En18
  input [18:0] Wgt_6_410, // sfix19_En18
  input [18:0] Wgt_6_411, // sfix19_En18
  input [18:0] Wgt_6_412, // sfix19_En18
  input [18:0] Wgt_6_413, // sfix19_En18
  input [18:0] Wgt_6_414, // sfix19_En18
  input [18:0] Wgt_6_415, // sfix19_En18
  input [18:0] Wgt_6_416, // sfix19_En18
  input [18:0] Wgt_6_417, // sfix19_En18
  input [18:0] Wgt_6_418, // sfix19_En18
  input [18:0] Wgt_6_419, // sfix19_En18
  input [18:0] Wgt_6_420, // sfix19_En18
  input [18:0] Wgt_6_421, // sfix19_En18
  input [18:0] Wgt_6_422, // sfix19_En18
  input [18:0] Wgt_6_423, // sfix19_En18
  input [18:0] Wgt_6_424, // sfix19_En18
  input [18:0] Wgt_6_425, // sfix19_En18
  input [18:0] Wgt_6_426, // sfix19_En18
  input [18:0] Wgt_6_427, // sfix19_En18
  input [18:0] Wgt_6_428, // sfix19_En18
  input [18:0] Wgt_6_429, // sfix19_En18
  input [18:0] Wgt_6_430, // sfix19_En18
  input [18:0] Wgt_6_431, // sfix19_En18
  input [18:0] Wgt_6_432, // sfix19_En18
  input [18:0] Wgt_6_433, // sfix19_En18
  input [18:0] Wgt_6_434, // sfix19_En18
  input [18:0] Wgt_6_435, // sfix19_En18
  input [18:0] Wgt_6_436, // sfix19_En18
  input [18:0] Wgt_6_437, // sfix19_En18
  input [18:0] Wgt_6_438, // sfix19_En18
  input [18:0] Wgt_6_439, // sfix19_En18
  input [18:0] Wgt_6_440, // sfix19_En18
  input [18:0] Wgt_6_441, // sfix19_En18
  input [18:0] Wgt_6_442, // sfix19_En18
  input [18:0] Wgt_6_443, // sfix19_En18
  input [18:0] Wgt_6_444, // sfix19_En18
  input [18:0] Wgt_6_445, // sfix19_En18
  input [18:0] Wgt_6_446, // sfix19_En18
  input [18:0] Wgt_6_447, // sfix19_En18
  input [18:0] Wgt_6_448, // sfix19_En18
  input [18:0] Wgt_6_449, // sfix19_En18
  input [18:0] Wgt_6_450, // sfix19_En18
  input [18:0] Wgt_6_451, // sfix19_En18
  input [18:0] Wgt_6_452, // sfix19_En18
  input [18:0] Wgt_6_453, // sfix19_En18
  input [18:0] Wgt_6_454, // sfix19_En18
  input [18:0] Wgt_6_455, // sfix19_En18
  input [18:0] Wgt_6_456, // sfix19_En18
  input [18:0] Wgt_6_457, // sfix19_En18
  input [18:0] Wgt_6_458, // sfix19_En18
  input [18:0] Wgt_6_459, // sfix19_En18
  input [18:0] Wgt_6_460, // sfix19_En18
  input [18:0] Wgt_6_461, // sfix19_En18
  input [18:0] Wgt_6_462, // sfix19_En18
  input [18:0] Wgt_6_463, // sfix19_En18
  input [18:0] Wgt_6_464, // sfix19_En18
  input [18:0] Wgt_6_465, // sfix19_En18
  input [18:0] Wgt_6_466, // sfix19_En18
  input [18:0] Wgt_6_467, // sfix19_En18
  input [18:0] Wgt_6_468, // sfix19_En18
  input [18:0] Wgt_6_469, // sfix19_En18
  input [18:0] Wgt_6_470, // sfix19_En18
  input [18:0] Wgt_6_471, // sfix19_En18
  input [18:0] Wgt_6_472, // sfix19_En18
  input [18:0] Wgt_6_473, // sfix19_En18
  input [18:0] Wgt_6_474, // sfix19_En18
  input [18:0] Wgt_6_475, // sfix19_En18
  input [18:0] Wgt_6_476, // sfix19_En18
  input [18:0] Wgt_6_477, // sfix19_En18
  input [18:0] Wgt_6_478, // sfix19_En18
  input [18:0] Wgt_6_479, // sfix19_En18
  input [18:0] Wgt_6_480, // sfix19_En18
  input [18:0] Wgt_6_481, // sfix19_En18
  input [18:0] Wgt_6_482, // sfix19_En18
  input [18:0] Wgt_6_483, // sfix19_En18
  input [18:0] Wgt_6_484, // sfix19_En18
  input [18:0] Wgt_6_485, // sfix19_En18
  input [18:0] Wgt_6_486, // sfix19_En18
  input [18:0] Wgt_6_487, // sfix19_En18
  input [18:0] Wgt_6_488, // sfix19_En18
  input [18:0] Wgt_6_489, // sfix19_En18
  input [18:0] Wgt_6_490, // sfix19_En18
  input [18:0] Wgt_6_491, // sfix19_En18
  input [18:0] Wgt_6_492, // sfix19_En18
  input [18:0] Wgt_6_493, // sfix19_En18
  input [18:0] Wgt_6_494, // sfix19_En18
  input [18:0] Wgt_6_495, // sfix19_En18
  input [18:0] Wgt_6_496, // sfix19_En18
  input [18:0] Wgt_6_497, // sfix19_En18
  input [18:0] Wgt_6_498, // sfix19_En18
  input [18:0] Wgt_6_499, // sfix19_En18
  input [18:0] Wgt_6_500, // sfix19_En18
  input [18:0] Wgt_6_501, // sfix19_En18
  input [18:0] Wgt_6_502, // sfix19_En18
  input [18:0] Wgt_6_503, // sfix19_En18
  input [18:0] Wgt_6_504, // sfix19_En18
  input [18:0] Wgt_6_505, // sfix19_En18
  input [18:0] Wgt_6_506, // sfix19_En18
  input [18:0] Wgt_6_507, // sfix19_En18
  input [18:0] Wgt_6_508, // sfix19_En18
  input [18:0] Wgt_6_509, // sfix19_En18
  input [18:0] Wgt_6_510, // sfix19_En18
  input [18:0] Wgt_6_511, // sfix19_En18
  input [18:0] Wgt_6_512, // sfix19_En18
  input [18:0] Wgt_6_513, // sfix19_En18
  input [18:0] Wgt_6_514, // sfix19_En18
  input [18:0] Wgt_6_515, // sfix19_En18
  input [18:0] Wgt_6_516, // sfix19_En18
  input [18:0] Wgt_6_517, // sfix19_En18
  input [18:0] Wgt_6_518, // sfix19_En18
  input [18:0] Wgt_6_519, // sfix19_En18
  input [18:0] Wgt_6_520, // sfix19_En18
  input [18:0] Wgt_6_521, // sfix19_En18
  input [18:0] Wgt_6_522, // sfix19_En18
  input [18:0] Wgt_6_523, // sfix19_En18
  input [18:0] Wgt_6_524, // sfix19_En18
  input [18:0] Wgt_6_525, // sfix19_En18
  input [18:0] Wgt_6_526, // sfix19_En18
  input [18:0] Wgt_6_527, // sfix19_En18
  input [18:0] Wgt_6_528, // sfix19_En18
  input [18:0] Wgt_6_529, // sfix19_En18
  input [18:0] Wgt_6_530, // sfix19_En18
  input [18:0] Wgt_6_531, // sfix19_En18
  input [18:0] Wgt_6_532, // sfix19_En18
  input [18:0] Wgt_6_533, // sfix19_En18
  input [18:0] Wgt_6_534, // sfix19_En18
  input [18:0] Wgt_6_535, // sfix19_En18
  input [18:0] Wgt_6_536, // sfix19_En18
  input [18:0] Wgt_6_537, // sfix19_En18
  input [18:0] Wgt_6_538, // sfix19_En18
  input [18:0] Wgt_6_539, // sfix19_En18
  input [18:0] Wgt_6_540, // sfix19_En18
  input [18:0] Wgt_6_541, // sfix19_En18
  input [18:0] Wgt_6_542, // sfix19_En18
  input [18:0] Wgt_6_543, // sfix19_En18
  input [18:0] Wgt_6_544, // sfix19_En18
  input [18:0] Wgt_6_545, // sfix19_En18
  input [18:0] Wgt_6_546, // sfix19_En18
  input [18:0] Wgt_6_547, // sfix19_En18
  input [18:0] Wgt_6_548, // sfix19_En18
  input [18:0] Wgt_6_549, // sfix19_En18
  input [18:0] Wgt_6_550, // sfix19_En18
  input [18:0] Wgt_6_551, // sfix19_En18
  input [18:0] Wgt_6_552, // sfix19_En18
  input [18:0] Wgt_6_553, // sfix19_En18
  input [18:0] Wgt_6_554, // sfix19_En18
  input [18:0] Wgt_6_555, // sfix19_En18
  input [18:0] Wgt_6_556, // sfix19_En18
  input [18:0] Wgt_6_557, // sfix19_En18
  input [18:0] Wgt_6_558, // sfix19_En18
  input [18:0] Wgt_6_559, // sfix19_En18
  input [18:0] Wgt_6_560, // sfix19_En18
  input [18:0] Wgt_6_561, // sfix19_En18
  input [18:0] Wgt_6_562, // sfix19_En18
  input [18:0] Wgt_6_563, // sfix19_En18
  input [18:0] Wgt_6_564, // sfix19_En18
  input [18:0] Wgt_6_565, // sfix19_En18
  input [18:0] Wgt_6_566, // sfix19_En18
  input [18:0] Wgt_6_567, // sfix19_En18
  input [18:0] Wgt_6_568, // sfix19_En18
  input [18:0] Wgt_6_569, // sfix19_En18
  input [18:0] Wgt_6_570, // sfix19_En18
  input [18:0] Wgt_6_571, // sfix19_En18
  input [18:0] Wgt_6_572, // sfix19_En18
  input [18:0] Wgt_6_573, // sfix19_En18
  input [18:0] Wgt_6_574, // sfix19_En18
  input [18:0] Wgt_6_575, // sfix19_En18
  input [18:0] Wgt_6_576, // sfix19_En18
  input [18:0] Wgt_6_577, // sfix19_En18
  input [18:0] Wgt_6_578, // sfix19_En18
  input [18:0] Wgt_6_579, // sfix19_En18
  input [18:0] Wgt_6_580, // sfix19_En18
  input [18:0] Wgt_6_581, // sfix19_En18
  input [18:0] Wgt_6_582, // sfix19_En18
  input [18:0] Wgt_6_583, // sfix19_En18
  input [18:0] Wgt_6_584, // sfix19_En18
  input [18:0] Wgt_6_585, // sfix19_En18
  input [18:0] Wgt_6_586, // sfix19_En18
  input [18:0] Wgt_6_587, // sfix19_En18
  input [18:0] Wgt_6_588, // sfix19_En18
  input [18:0] Wgt_6_589, // sfix19_En18
  input [18:0] Wgt_6_590, // sfix19_En18
  input [18:0] Wgt_6_591, // sfix19_En18
  input [18:0] Wgt_6_592, // sfix19_En18
  input [18:0] Wgt_6_593, // sfix19_En18
  input [18:0] Wgt_6_594, // sfix19_En18
  input [18:0] Wgt_6_595, // sfix19_En18
  input [18:0] Wgt_6_596, // sfix19_En18
  input [18:0] Wgt_6_597, // sfix19_En18
  input [18:0] Wgt_6_598, // sfix19_En18
  input [18:0] Wgt_6_599, // sfix19_En18
  input [18:0] Wgt_6_600, // sfix19_En18
  input [18:0] Wgt_6_601, // sfix19_En18
  input [18:0] Wgt_6_602, // sfix19_En18
  input [18:0] Wgt_6_603, // sfix19_En18
  input [18:0] Wgt_6_604, // sfix19_En18
  input [18:0] Wgt_6_605, // sfix19_En18
  input [18:0] Wgt_6_606, // sfix19_En18
  input [18:0] Wgt_6_607, // sfix19_En18
  input [18:0] Wgt_6_608, // sfix19_En18
  input [18:0] Wgt_6_609, // sfix19_En18
  input [18:0] Wgt_6_610, // sfix19_En18
  input [18:0] Wgt_6_611, // sfix19_En18
  input [18:0] Wgt_6_612, // sfix19_En18
  input [18:0] Wgt_6_613, // sfix19_En18
  input [18:0] Wgt_6_614, // sfix19_En18
  input [18:0] Wgt_6_615, // sfix19_En18
  input [18:0] Wgt_6_616, // sfix19_En18
  input [18:0] Wgt_6_617, // sfix19_En18
  input [18:0] Wgt_6_618, // sfix19_En18
  input [18:0] Wgt_6_619, // sfix19_En18
  input [18:0] Wgt_6_620, // sfix19_En18
  input [18:0] Wgt_6_621, // sfix19_En18
  input [18:0] Wgt_6_622, // sfix19_En18
  input [18:0] Wgt_6_623, // sfix19_En18
  input [18:0] Wgt_6_624, // sfix19_En18
  input [18:0] Wgt_6_625, // sfix19_En18
  input [18:0] Wgt_6_626, // sfix19_En18
  input [18:0] Wgt_6_627, // sfix19_En18
  input [18:0] Wgt_6_628, // sfix19_En18
  input [18:0] Wgt_6_629, // sfix19_En18
  input [18:0] Wgt_6_630, // sfix19_En18
  input [18:0] Wgt_6_631, // sfix19_En18
  input [18:0] Wgt_6_632, // sfix19_En18
  input [18:0] Wgt_6_633, // sfix19_En18
  input [18:0] Wgt_6_634, // sfix19_En18
  input [18:0] Wgt_6_635, // sfix19_En18
  input [18:0] Wgt_6_636, // sfix19_En18
  input [18:0] Wgt_6_637, // sfix19_En18
  input [18:0] Wgt_6_638, // sfix19_En18
  input [18:0] Wgt_6_639, // sfix19_En18
  input [18:0] Wgt_6_640, // sfix19_En18
  input [18:0] Wgt_6_641, // sfix19_En18
  input [18:0] Wgt_6_642, // sfix19_En18
  input [18:0] Wgt_6_643, // sfix19_En18
  input [18:0] Wgt_6_644, // sfix19_En18
  input [18:0] Wgt_6_645, // sfix19_En18
  input [18:0] Wgt_6_646, // sfix19_En18
  input [18:0] Wgt_6_647, // sfix19_En18
  input [18:0] Wgt_6_648, // sfix19_En18
  input [18:0] Wgt_6_649, // sfix19_En18
  input [18:0] Wgt_6_650, // sfix19_En18
  input [18:0] Wgt_6_651, // sfix19_En18
  input [18:0] Wgt_6_652, // sfix19_En18
  input [18:0] Wgt_6_653, // sfix19_En18
  input [18:0] Wgt_6_654, // sfix19_En18
  input [18:0] Wgt_6_655, // sfix19_En18
  input [18:0] Wgt_6_656, // sfix19_En18
  input [18:0] Wgt_6_657, // sfix19_En18
  input [18:0] Wgt_6_658, // sfix19_En18
  input [18:0] Wgt_6_659, // sfix19_En18
  input [18:0] Wgt_6_660, // sfix19_En18
  input [18:0] Wgt_6_661, // sfix19_En18
  input [18:0] Wgt_6_662, // sfix19_En18
  input [18:0] Wgt_6_663, // sfix19_En18
  input [18:0] Wgt_6_664, // sfix19_En18
  input [18:0] Wgt_6_665, // sfix19_En18
  input [18:0] Wgt_6_666, // sfix19_En18
  input [18:0] Wgt_6_667, // sfix19_En18
  input [18:0] Wgt_6_668, // sfix19_En18
  input [18:0] Wgt_6_669, // sfix19_En18
  input [18:0] Wgt_6_670, // sfix19_En18
  input [18:0] Wgt_6_671, // sfix19_En18
  input [18:0] Wgt_6_672, // sfix19_En18
  input [18:0] Wgt_6_673, // sfix19_En18
  input [18:0] Wgt_6_674, // sfix19_En18
  input [18:0] Wgt_6_675, // sfix19_En18
  input [18:0] Wgt_6_676, // sfix19_En18
  input [18:0] Wgt_6_677, // sfix19_En18
  input [18:0] Wgt_6_678, // sfix19_En18
  input [18:0] Wgt_6_679, // sfix19_En18
  input [18:0] Wgt_6_680, // sfix19_En18
  input [18:0] Wgt_6_681, // sfix19_En18
  input [18:0] Wgt_6_682, // sfix19_En18
  input [18:0] Wgt_6_683, // sfix19_En18
  input [18:0] Wgt_6_684, // sfix19_En18
  input [18:0] Wgt_6_685, // sfix19_En18
  input [18:0] Wgt_6_686, // sfix19_En18
  input [18:0] Wgt_6_687, // sfix19_En18
  input [18:0] Wgt_6_688, // sfix19_En18
  input [18:0] Wgt_6_689, // sfix19_En18
  input [18:0] Wgt_6_690, // sfix19_En18
  input [18:0] Wgt_6_691, // sfix19_En18
  input [18:0] Wgt_6_692, // sfix19_En18
  input [18:0] Wgt_6_693, // sfix19_En18
  input [18:0] Wgt_6_694, // sfix19_En18
  input [18:0] Wgt_6_695, // sfix19_En18
  input [18:0] Wgt_6_696, // sfix19_En18
  input [18:0] Wgt_6_697, // sfix19_En18
  input [18:0] Wgt_6_698, // sfix19_En18
  input [18:0] Wgt_6_699, // sfix19_En18
  input [18:0] Wgt_6_700, // sfix19_En18
  input [18:0] Wgt_6_701, // sfix19_En18
  input [18:0] Wgt_6_702, // sfix19_En18
  input [18:0] Wgt_6_703, // sfix19_En18
  input [18:0] Wgt_6_704, // sfix19_En18
  input [18:0] Wgt_6_705, // sfix19_En18
  input [18:0] Wgt_6_706, // sfix19_En18
  input [18:0] Wgt_6_707, // sfix19_En18
  input [18:0] Wgt_6_708, // sfix19_En18
  input [18:0] Wgt_6_709, // sfix19_En18
  input [18:0] Wgt_6_710, // sfix19_En18
  input [18:0] Wgt_6_711, // sfix19_En18
  input [18:0] Wgt_6_712, // sfix19_En18
  input [18:0] Wgt_6_713, // sfix19_En18
  input [18:0] Wgt_6_714, // sfix19_En18
  input [18:0] Wgt_6_715, // sfix19_En18
  input [18:0] Wgt_6_716, // sfix19_En18
  input [18:0] Wgt_6_717, // sfix19_En18
  input [18:0] Wgt_6_718, // sfix19_En18
  input [18:0] Wgt_6_719, // sfix19_En18
  input [18:0] Wgt_6_720, // sfix19_En18
  input [18:0] Wgt_6_721, // sfix19_En18
  input [18:0] Wgt_6_722, // sfix19_En18
  input [18:0] Wgt_6_723, // sfix19_En18
  input [18:0] Wgt_6_724, // sfix19_En18
  input [18:0] Wgt_6_725, // sfix19_En18
  input [18:0] Wgt_6_726, // sfix19_En18
  input [18:0] Wgt_6_727, // sfix19_En18
  input [18:0] Wgt_6_728, // sfix19_En18
  input [18:0] Wgt_6_729, // sfix19_En18
  input [18:0] Wgt_6_730, // sfix19_En18
  input [18:0] Wgt_6_731, // sfix19_En18
  input [18:0] Wgt_6_732, // sfix19_En18
  input [18:0] Wgt_6_733, // sfix19_En18
  input [18:0] Wgt_6_734, // sfix19_En18
  input [18:0] Wgt_6_735, // sfix19_En18
  input [18:0] Wgt_6_736, // sfix19_En18
  input [18:0] Wgt_6_737, // sfix19_En18
  input [18:0] Wgt_6_738, // sfix19_En18
  input [18:0] Wgt_6_739, // sfix19_En18
  input [18:0] Wgt_6_740, // sfix19_En18
  input [18:0] Wgt_6_741, // sfix19_En18
  input [18:0] Wgt_6_742, // sfix19_En18
  input [18:0] Wgt_6_743, // sfix19_En18
  input [18:0] Wgt_6_744, // sfix19_En18
  input [18:0] Wgt_6_745, // sfix19_En18
  input [18:0] Wgt_6_746, // sfix19_En18
  input [18:0] Wgt_6_747, // sfix19_En18
  input [18:0] Wgt_6_748, // sfix19_En18
  input [18:0] Wgt_6_749, // sfix19_En18
  input [18:0] Wgt_6_750, // sfix19_En18
  input [18:0] Wgt_6_751, // sfix19_En18
  input [18:0] Wgt_6_752, // sfix19_En18
  input [18:0] Wgt_6_753, // sfix19_En18
  input [18:0] Wgt_6_754, // sfix19_En18
  input [18:0] Wgt_6_755, // sfix19_En18
  input [18:0] Wgt_6_756, // sfix19_En18
  input [18:0] Wgt_6_757, // sfix19_En18
  input [18:0] Wgt_6_758, // sfix19_En18
  input [18:0] Wgt_6_759, // sfix19_En18
  input [18:0] Wgt_6_760, // sfix19_En18
  input [18:0] Wgt_6_761, // sfix19_En18
  input [18:0] Wgt_6_762, // sfix19_En18
  input [18:0] Wgt_6_763, // sfix19_En18
  input [18:0] Wgt_6_764, // sfix19_En18
  input [18:0] Wgt_6_765, // sfix19_En18
  input [18:0] Wgt_6_766, // sfix19_En18
  input [18:0] Wgt_6_767, // sfix19_En18
  input [18:0] Wgt_6_768, // sfix19_En18
  input [18:0] Wgt_6_769, // sfix19_En18
  input [18:0] Wgt_6_770, // sfix19_En18
  input [18:0] Wgt_6_771, // sfix19_En18
  input [18:0] Wgt_6_772, // sfix19_En18
  input [18:0] Wgt_6_773, // sfix19_En18
  input [18:0] Wgt_6_774, // sfix19_En18
  input [18:0] Wgt_6_775, // sfix19_En18
  input [18:0] Wgt_6_776, // sfix19_En18
  input [18:0] Wgt_6_777, // sfix19_En18
  input [18:0] Wgt_6_778, // sfix19_En18
  input [18:0] Wgt_6_779, // sfix19_En18
  input [18:0] Wgt_6_780, // sfix19_En18
  input [18:0] Wgt_6_781, // sfix19_En18
  input [18:0] Wgt_6_782, // sfix19_En18
  input [18:0] Wgt_6_783, // sfix19_En18
  input [18:0] Wgt_6_784, // sfix19_En18
  input [18:0] Wgt_7_0, // sfix19_En18
  input [18:0] Wgt_7_1, // sfix19_En18
  input [18:0] Wgt_7_2, // sfix19_En18
  input [18:0] Wgt_7_3, // sfix19_En18
  input [18:0] Wgt_7_4, // sfix19_En18
  input [18:0] Wgt_7_5, // sfix19_En18
  input [18:0] Wgt_7_6, // sfix19_En18
  input [18:0] Wgt_7_7, // sfix19_En18
  input [18:0] Wgt_7_8, // sfix19_En18
  input [18:0] Wgt_7_9, // sfix19_En18
  input [18:0] Wgt_7_10, // sfix19_En18
  input [18:0] Wgt_7_11, // sfix19_En18
  input [18:0] Wgt_7_12, // sfix19_En18
  input [18:0] Wgt_7_13, // sfix19_En18
  input [18:0] Wgt_7_14, // sfix19_En18
  input [18:0] Wgt_7_15, // sfix19_En18
  input [18:0] Wgt_7_16, // sfix19_En18
  input [18:0] Wgt_7_17, // sfix19_En18
  input [18:0] Wgt_7_18, // sfix19_En18
  input [18:0] Wgt_7_19, // sfix19_En18
  input [18:0] Wgt_7_20, // sfix19_En18
  input [18:0] Wgt_7_21, // sfix19_En18
  input [18:0] Wgt_7_22, // sfix19_En18
  input [18:0] Wgt_7_23, // sfix19_En18
  input [18:0] Wgt_7_24, // sfix19_En18
  input [18:0] Wgt_7_25, // sfix19_En18
  input [18:0] Wgt_7_26, // sfix19_En18
  input [18:0] Wgt_7_27, // sfix19_En18
  input [18:0] Wgt_7_28, // sfix19_En18
  input [18:0] Wgt_7_29, // sfix19_En18
  input [18:0] Wgt_7_30, // sfix19_En18
  input [18:0] Wgt_7_31, // sfix19_En18
  input [18:0] Wgt_7_32, // sfix19_En18
  input [18:0] Wgt_7_33, // sfix19_En18
  input [18:0] Wgt_7_34, // sfix19_En18
  input [18:0] Wgt_7_35, // sfix19_En18
  input [18:0] Wgt_7_36, // sfix19_En18
  input [18:0] Wgt_7_37, // sfix19_En18
  input [18:0] Wgt_7_38, // sfix19_En18
  input [18:0] Wgt_7_39, // sfix19_En18
  input [18:0] Wgt_7_40, // sfix19_En18
  input [18:0] Wgt_7_41, // sfix19_En18
  input [18:0] Wgt_7_42, // sfix19_En18
  input [18:0] Wgt_7_43, // sfix19_En18
  input [18:0] Wgt_7_44, // sfix19_En18
  input [18:0] Wgt_7_45, // sfix19_En18
  input [18:0] Wgt_7_46, // sfix19_En18
  input [18:0] Wgt_7_47, // sfix19_En18
  input [18:0] Wgt_7_48, // sfix19_En18
  input [18:0] Wgt_7_49, // sfix19_En18
  input [18:0] Wgt_7_50, // sfix19_En18
  input [18:0] Wgt_7_51, // sfix19_En18
  input [18:0] Wgt_7_52, // sfix19_En18
  input [18:0] Wgt_7_53, // sfix19_En18
  input [18:0] Wgt_7_54, // sfix19_En18
  input [18:0] Wgt_7_55, // sfix19_En18
  input [18:0] Wgt_7_56, // sfix19_En18
  input [18:0] Wgt_7_57, // sfix19_En18
  input [18:0] Wgt_7_58, // sfix19_En18
  input [18:0] Wgt_7_59, // sfix19_En18
  input [18:0] Wgt_7_60, // sfix19_En18
  input [18:0] Wgt_7_61, // sfix19_En18
  input [18:0] Wgt_7_62, // sfix19_En18
  input [18:0] Wgt_7_63, // sfix19_En18
  input [18:0] Wgt_7_64, // sfix19_En18
  input [18:0] Wgt_7_65, // sfix19_En18
  input [18:0] Wgt_7_66, // sfix19_En18
  input [18:0] Wgt_7_67, // sfix19_En18
  input [18:0] Wgt_7_68, // sfix19_En18
  input [18:0] Wgt_7_69, // sfix19_En18
  input [18:0] Wgt_7_70, // sfix19_En18
  input [18:0] Wgt_7_71, // sfix19_En18
  input [18:0] Wgt_7_72, // sfix19_En18
  input [18:0] Wgt_7_73, // sfix19_En18
  input [18:0] Wgt_7_74, // sfix19_En18
  input [18:0] Wgt_7_75, // sfix19_En18
  input [18:0] Wgt_7_76, // sfix19_En18
  input [18:0] Wgt_7_77, // sfix19_En18
  input [18:0] Wgt_7_78, // sfix19_En18
  input [18:0] Wgt_7_79, // sfix19_En18
  input [18:0] Wgt_7_80, // sfix19_En18
  input [18:0] Wgt_7_81, // sfix19_En18
  input [18:0] Wgt_7_82, // sfix19_En18
  input [18:0] Wgt_7_83, // sfix19_En18
  input [18:0] Wgt_7_84, // sfix19_En18
  input [18:0] Wgt_7_85, // sfix19_En18
  input [18:0] Wgt_7_86, // sfix19_En18
  input [18:0] Wgt_7_87, // sfix19_En18
  input [18:0] Wgt_7_88, // sfix19_En18
  input [18:0] Wgt_7_89, // sfix19_En18
  input [18:0] Wgt_7_90, // sfix19_En18
  input [18:0] Wgt_7_91, // sfix19_En18
  input [18:0] Wgt_7_92, // sfix19_En18
  input [18:0] Wgt_7_93, // sfix19_En18
  input [18:0] Wgt_7_94, // sfix19_En18
  input [18:0] Wgt_7_95, // sfix19_En18
  input [18:0] Wgt_7_96, // sfix19_En18
  input [18:0] Wgt_7_97, // sfix19_En18
  input [18:0] Wgt_7_98, // sfix19_En18
  input [18:0] Wgt_7_99, // sfix19_En18
  input [18:0] Wgt_7_100, // sfix19_En18
  input [18:0] Wgt_7_101, // sfix19_En18
  input [18:0] Wgt_7_102, // sfix19_En18
  input [18:0] Wgt_7_103, // sfix19_En18
  input [18:0] Wgt_7_104, // sfix19_En18
  input [18:0] Wgt_7_105, // sfix19_En18
  input [18:0] Wgt_7_106, // sfix19_En18
  input [18:0] Wgt_7_107, // sfix19_En18
  input [18:0] Wgt_7_108, // sfix19_En18
  input [18:0] Wgt_7_109, // sfix19_En18
  input [18:0] Wgt_7_110, // sfix19_En18
  input [18:0] Wgt_7_111, // sfix19_En18
  input [18:0] Wgt_7_112, // sfix19_En18
  input [18:0] Wgt_7_113, // sfix19_En18
  input [18:0] Wgt_7_114, // sfix19_En18
  input [18:0] Wgt_7_115, // sfix19_En18
  input [18:0] Wgt_7_116, // sfix19_En18
  input [18:0] Wgt_7_117, // sfix19_En18
  input [18:0] Wgt_7_118, // sfix19_En18
  input [18:0] Wgt_7_119, // sfix19_En18
  input [18:0] Wgt_7_120, // sfix19_En18
  input [18:0] Wgt_7_121, // sfix19_En18
  input [18:0] Wgt_7_122, // sfix19_En18
  input [18:0] Wgt_7_123, // sfix19_En18
  input [18:0] Wgt_7_124, // sfix19_En18
  input [18:0] Wgt_7_125, // sfix19_En18
  input [18:0] Wgt_7_126, // sfix19_En18
  input [18:0] Wgt_7_127, // sfix19_En18
  input [18:0] Wgt_7_128, // sfix19_En18
  input [18:0] Wgt_7_129, // sfix19_En18
  input [18:0] Wgt_7_130, // sfix19_En18
  input [18:0] Wgt_7_131, // sfix19_En18
  input [18:0] Wgt_7_132, // sfix19_En18
  input [18:0] Wgt_7_133, // sfix19_En18
  input [18:0] Wgt_7_134, // sfix19_En18
  input [18:0] Wgt_7_135, // sfix19_En18
  input [18:0] Wgt_7_136, // sfix19_En18
  input [18:0] Wgt_7_137, // sfix19_En18
  input [18:0] Wgt_7_138, // sfix19_En18
  input [18:0] Wgt_7_139, // sfix19_En18
  input [18:0] Wgt_7_140, // sfix19_En18
  input [18:0] Wgt_7_141, // sfix19_En18
  input [18:0] Wgt_7_142, // sfix19_En18
  input [18:0] Wgt_7_143, // sfix19_En18
  input [18:0] Wgt_7_144, // sfix19_En18
  input [18:0] Wgt_7_145, // sfix19_En18
  input [18:0] Wgt_7_146, // sfix19_En18
  input [18:0] Wgt_7_147, // sfix19_En18
  input [18:0] Wgt_7_148, // sfix19_En18
  input [18:0] Wgt_7_149, // sfix19_En18
  input [18:0] Wgt_7_150, // sfix19_En18
  input [18:0] Wgt_7_151, // sfix19_En18
  input [18:0] Wgt_7_152, // sfix19_En18
  input [18:0] Wgt_7_153, // sfix19_En18
  input [18:0] Wgt_7_154, // sfix19_En18
  input [18:0] Wgt_7_155, // sfix19_En18
  input [18:0] Wgt_7_156, // sfix19_En18
  input [18:0] Wgt_7_157, // sfix19_En18
  input [18:0] Wgt_7_158, // sfix19_En18
  input [18:0] Wgt_7_159, // sfix19_En18
  input [18:0] Wgt_7_160, // sfix19_En18
  input [18:0] Wgt_7_161, // sfix19_En18
  input [18:0] Wgt_7_162, // sfix19_En18
  input [18:0] Wgt_7_163, // sfix19_En18
  input [18:0] Wgt_7_164, // sfix19_En18
  input [18:0] Wgt_7_165, // sfix19_En18
  input [18:0] Wgt_7_166, // sfix19_En18
  input [18:0] Wgt_7_167, // sfix19_En18
  input [18:0] Wgt_7_168, // sfix19_En18
  input [18:0] Wgt_7_169, // sfix19_En18
  input [18:0] Wgt_7_170, // sfix19_En18
  input [18:0] Wgt_7_171, // sfix19_En18
  input [18:0] Wgt_7_172, // sfix19_En18
  input [18:0] Wgt_7_173, // sfix19_En18
  input [18:0] Wgt_7_174, // sfix19_En18
  input [18:0] Wgt_7_175, // sfix19_En18
  input [18:0] Wgt_7_176, // sfix19_En18
  input [18:0] Wgt_7_177, // sfix19_En18
  input [18:0] Wgt_7_178, // sfix19_En18
  input [18:0] Wgt_7_179, // sfix19_En18
  input [18:0] Wgt_7_180, // sfix19_En18
  input [18:0] Wgt_7_181, // sfix19_En18
  input [18:0] Wgt_7_182, // sfix19_En18
  input [18:0] Wgt_7_183, // sfix19_En18
  input [18:0] Wgt_7_184, // sfix19_En18
  input [18:0] Wgt_7_185, // sfix19_En18
  input [18:0] Wgt_7_186, // sfix19_En18
  input [18:0] Wgt_7_187, // sfix19_En18
  input [18:0] Wgt_7_188, // sfix19_En18
  input [18:0] Wgt_7_189, // sfix19_En18
  input [18:0] Wgt_7_190, // sfix19_En18
  input [18:0] Wgt_7_191, // sfix19_En18
  input [18:0] Wgt_7_192, // sfix19_En18
  input [18:0] Wgt_7_193, // sfix19_En18
  input [18:0] Wgt_7_194, // sfix19_En18
  input [18:0] Wgt_7_195, // sfix19_En18
  input [18:0] Wgt_7_196, // sfix19_En18
  input [18:0] Wgt_7_197, // sfix19_En18
  input [18:0] Wgt_7_198, // sfix19_En18
  input [18:0] Wgt_7_199, // sfix19_En18
  input [18:0] Wgt_7_200, // sfix19_En18
  input [18:0] Wgt_7_201, // sfix19_En18
  input [18:0] Wgt_7_202, // sfix19_En18
  input [18:0] Wgt_7_203, // sfix19_En18
  input [18:0] Wgt_7_204, // sfix19_En18
  input [18:0] Wgt_7_205, // sfix19_En18
  input [18:0] Wgt_7_206, // sfix19_En18
  input [18:0] Wgt_7_207, // sfix19_En18
  input [18:0] Wgt_7_208, // sfix19_En18
  input [18:0] Wgt_7_209, // sfix19_En18
  input [18:0] Wgt_7_210, // sfix19_En18
  input [18:0] Wgt_7_211, // sfix19_En18
  input [18:0] Wgt_7_212, // sfix19_En18
  input [18:0] Wgt_7_213, // sfix19_En18
  input [18:0] Wgt_7_214, // sfix19_En18
  input [18:0] Wgt_7_215, // sfix19_En18
  input [18:0] Wgt_7_216, // sfix19_En18
  input [18:0] Wgt_7_217, // sfix19_En18
  input [18:0] Wgt_7_218, // sfix19_En18
  input [18:0] Wgt_7_219, // sfix19_En18
  input [18:0] Wgt_7_220, // sfix19_En18
  input [18:0] Wgt_7_221, // sfix19_En18
  input [18:0] Wgt_7_222, // sfix19_En18
  input [18:0] Wgt_7_223, // sfix19_En18
  input [18:0] Wgt_7_224, // sfix19_En18
  input [18:0] Wgt_7_225, // sfix19_En18
  input [18:0] Wgt_7_226, // sfix19_En18
  input [18:0] Wgt_7_227, // sfix19_En18
  input [18:0] Wgt_7_228, // sfix19_En18
  input [18:0] Wgt_7_229, // sfix19_En18
  input [18:0] Wgt_7_230, // sfix19_En18
  input [18:0] Wgt_7_231, // sfix19_En18
  input [18:0] Wgt_7_232, // sfix19_En18
  input [18:0] Wgt_7_233, // sfix19_En18
  input [18:0] Wgt_7_234, // sfix19_En18
  input [18:0] Wgt_7_235, // sfix19_En18
  input [18:0] Wgt_7_236, // sfix19_En18
  input [18:0] Wgt_7_237, // sfix19_En18
  input [18:0] Wgt_7_238, // sfix19_En18
  input [18:0] Wgt_7_239, // sfix19_En18
  input [18:0] Wgt_7_240, // sfix19_En18
  input [18:0] Wgt_7_241, // sfix19_En18
  input [18:0] Wgt_7_242, // sfix19_En18
  input [18:0] Wgt_7_243, // sfix19_En18
  input [18:0] Wgt_7_244, // sfix19_En18
  input [18:0] Wgt_7_245, // sfix19_En18
  input [18:0] Wgt_7_246, // sfix19_En18
  input [18:0] Wgt_7_247, // sfix19_En18
  input [18:0] Wgt_7_248, // sfix19_En18
  input [18:0] Wgt_7_249, // sfix19_En18
  input [18:0] Wgt_7_250, // sfix19_En18
  input [18:0] Wgt_7_251, // sfix19_En18
  input [18:0] Wgt_7_252, // sfix19_En18
  input [18:0] Wgt_7_253, // sfix19_En18
  input [18:0] Wgt_7_254, // sfix19_En18
  input [18:0] Wgt_7_255, // sfix19_En18
  input [18:0] Wgt_7_256, // sfix19_En18
  input [18:0] Wgt_7_257, // sfix19_En18
  input [18:0] Wgt_7_258, // sfix19_En18
  input [18:0] Wgt_7_259, // sfix19_En18
  input [18:0] Wgt_7_260, // sfix19_En18
  input [18:0] Wgt_7_261, // sfix19_En18
  input [18:0] Wgt_7_262, // sfix19_En18
  input [18:0] Wgt_7_263, // sfix19_En18
  input [18:0] Wgt_7_264, // sfix19_En18
  input [18:0] Wgt_7_265, // sfix19_En18
  input [18:0] Wgt_7_266, // sfix19_En18
  input [18:0] Wgt_7_267, // sfix19_En18
  input [18:0] Wgt_7_268, // sfix19_En18
  input [18:0] Wgt_7_269, // sfix19_En18
  input [18:0] Wgt_7_270, // sfix19_En18
  input [18:0] Wgt_7_271, // sfix19_En18
  input [18:0] Wgt_7_272, // sfix19_En18
  input [18:0] Wgt_7_273, // sfix19_En18
  input [18:0] Wgt_7_274, // sfix19_En18
  input [18:0] Wgt_7_275, // sfix19_En18
  input [18:0] Wgt_7_276, // sfix19_En18
  input [18:0] Wgt_7_277, // sfix19_En18
  input [18:0] Wgt_7_278, // sfix19_En18
  input [18:0] Wgt_7_279, // sfix19_En18
  input [18:0] Wgt_7_280, // sfix19_En18
  input [18:0] Wgt_7_281, // sfix19_En18
  input [18:0] Wgt_7_282, // sfix19_En18
  input [18:0] Wgt_7_283, // sfix19_En18
  input [18:0] Wgt_7_284, // sfix19_En18
  input [18:0] Wgt_7_285, // sfix19_En18
  input [18:0] Wgt_7_286, // sfix19_En18
  input [18:0] Wgt_7_287, // sfix19_En18
  input [18:0] Wgt_7_288, // sfix19_En18
  input [18:0] Wgt_7_289, // sfix19_En18
  input [18:0] Wgt_7_290, // sfix19_En18
  input [18:0] Wgt_7_291, // sfix19_En18
  input [18:0] Wgt_7_292, // sfix19_En18
  input [18:0] Wgt_7_293, // sfix19_En18
  input [18:0] Wgt_7_294, // sfix19_En18
  input [18:0] Wgt_7_295, // sfix19_En18
  input [18:0] Wgt_7_296, // sfix19_En18
  input [18:0] Wgt_7_297, // sfix19_En18
  input [18:0] Wgt_7_298, // sfix19_En18
  input [18:0] Wgt_7_299, // sfix19_En18
  input [18:0] Wgt_7_300, // sfix19_En18
  input [18:0] Wgt_7_301, // sfix19_En18
  input [18:0] Wgt_7_302, // sfix19_En18
  input [18:0] Wgt_7_303, // sfix19_En18
  input [18:0] Wgt_7_304, // sfix19_En18
  input [18:0] Wgt_7_305, // sfix19_En18
  input [18:0] Wgt_7_306, // sfix19_En18
  input [18:0] Wgt_7_307, // sfix19_En18
  input [18:0] Wgt_7_308, // sfix19_En18
  input [18:0] Wgt_7_309, // sfix19_En18
  input [18:0] Wgt_7_310, // sfix19_En18
  input [18:0] Wgt_7_311, // sfix19_En18
  input [18:0] Wgt_7_312, // sfix19_En18
  input [18:0] Wgt_7_313, // sfix19_En18
  input [18:0] Wgt_7_314, // sfix19_En18
  input [18:0] Wgt_7_315, // sfix19_En18
  input [18:0] Wgt_7_316, // sfix19_En18
  input [18:0] Wgt_7_317, // sfix19_En18
  input [18:0] Wgt_7_318, // sfix19_En18
  input [18:0] Wgt_7_319, // sfix19_En18
  input [18:0] Wgt_7_320, // sfix19_En18
  input [18:0] Wgt_7_321, // sfix19_En18
  input [18:0] Wgt_7_322, // sfix19_En18
  input [18:0] Wgt_7_323, // sfix19_En18
  input [18:0] Wgt_7_324, // sfix19_En18
  input [18:0] Wgt_7_325, // sfix19_En18
  input [18:0] Wgt_7_326, // sfix19_En18
  input [18:0] Wgt_7_327, // sfix19_En18
  input [18:0] Wgt_7_328, // sfix19_En18
  input [18:0] Wgt_7_329, // sfix19_En18
  input [18:0] Wgt_7_330, // sfix19_En18
  input [18:0] Wgt_7_331, // sfix19_En18
  input [18:0] Wgt_7_332, // sfix19_En18
  input [18:0] Wgt_7_333, // sfix19_En18
  input [18:0] Wgt_7_334, // sfix19_En18
  input [18:0] Wgt_7_335, // sfix19_En18
  input [18:0] Wgt_7_336, // sfix19_En18
  input [18:0] Wgt_7_337, // sfix19_En18
  input [18:0] Wgt_7_338, // sfix19_En18
  input [18:0] Wgt_7_339, // sfix19_En18
  input [18:0] Wgt_7_340, // sfix19_En18
  input [18:0] Wgt_7_341, // sfix19_En18
  input [18:0] Wgt_7_342, // sfix19_En18
  input [18:0] Wgt_7_343, // sfix19_En18
  input [18:0] Wgt_7_344, // sfix19_En18
  input [18:0] Wgt_7_345, // sfix19_En18
  input [18:0] Wgt_7_346, // sfix19_En18
  input [18:0] Wgt_7_347, // sfix19_En18
  input [18:0] Wgt_7_348, // sfix19_En18
  input [18:0] Wgt_7_349, // sfix19_En18
  input [18:0] Wgt_7_350, // sfix19_En18
  input [18:0] Wgt_7_351, // sfix19_En18
  input [18:0] Wgt_7_352, // sfix19_En18
  input [18:0] Wgt_7_353, // sfix19_En18
  input [18:0] Wgt_7_354, // sfix19_En18
  input [18:0] Wgt_7_355, // sfix19_En18
  input [18:0] Wgt_7_356, // sfix19_En18
  input [18:0] Wgt_7_357, // sfix19_En18
  input [18:0] Wgt_7_358, // sfix19_En18
  input [18:0] Wgt_7_359, // sfix19_En18
  input [18:0] Wgt_7_360, // sfix19_En18
  input [18:0] Wgt_7_361, // sfix19_En18
  input [18:0] Wgt_7_362, // sfix19_En18
  input [18:0] Wgt_7_363, // sfix19_En18
  input [18:0] Wgt_7_364, // sfix19_En18
  input [18:0] Wgt_7_365, // sfix19_En18
  input [18:0] Wgt_7_366, // sfix19_En18
  input [18:0] Wgt_7_367, // sfix19_En18
  input [18:0] Wgt_7_368, // sfix19_En18
  input [18:0] Wgt_7_369, // sfix19_En18
  input [18:0] Wgt_7_370, // sfix19_En18
  input [18:0] Wgt_7_371, // sfix19_En18
  input [18:0] Wgt_7_372, // sfix19_En18
  input [18:0] Wgt_7_373, // sfix19_En18
  input [18:0] Wgt_7_374, // sfix19_En18
  input [18:0] Wgt_7_375, // sfix19_En18
  input [18:0] Wgt_7_376, // sfix19_En18
  input [18:0] Wgt_7_377, // sfix19_En18
  input [18:0] Wgt_7_378, // sfix19_En18
  input [18:0] Wgt_7_379, // sfix19_En18
  input [18:0] Wgt_7_380, // sfix19_En18
  input [18:0] Wgt_7_381, // sfix19_En18
  input [18:0] Wgt_7_382, // sfix19_En18
  input [18:0] Wgt_7_383, // sfix19_En18
  input [18:0] Wgt_7_384, // sfix19_En18
  input [18:0] Wgt_7_385, // sfix19_En18
  input [18:0] Wgt_7_386, // sfix19_En18
  input [18:0] Wgt_7_387, // sfix19_En18
  input [18:0] Wgt_7_388, // sfix19_En18
  input [18:0] Wgt_7_389, // sfix19_En18
  input [18:0] Wgt_7_390, // sfix19_En18
  input [18:0] Wgt_7_391, // sfix19_En18
  input [18:0] Wgt_7_392, // sfix19_En18
  input [18:0] Wgt_7_393, // sfix19_En18
  input [18:0] Wgt_7_394, // sfix19_En18
  input [18:0] Wgt_7_395, // sfix19_En18
  input [18:0] Wgt_7_396, // sfix19_En18
  input [18:0] Wgt_7_397, // sfix19_En18
  input [18:0] Wgt_7_398, // sfix19_En18
  input [18:0] Wgt_7_399, // sfix19_En18
  input [18:0] Wgt_7_400, // sfix19_En18
  input [18:0] Wgt_7_401, // sfix19_En18
  input [18:0] Wgt_7_402, // sfix19_En18
  input [18:0] Wgt_7_403, // sfix19_En18
  input [18:0] Wgt_7_404, // sfix19_En18
  input [18:0] Wgt_7_405, // sfix19_En18
  input [18:0] Wgt_7_406, // sfix19_En18
  input [18:0] Wgt_7_407, // sfix19_En18
  input [18:0] Wgt_7_408, // sfix19_En18
  input [18:0] Wgt_7_409, // sfix19_En18
  input [18:0] Wgt_7_410, // sfix19_En18
  input [18:0] Wgt_7_411, // sfix19_En18
  input [18:0] Wgt_7_412, // sfix19_En18
  input [18:0] Wgt_7_413, // sfix19_En18
  input [18:0] Wgt_7_414, // sfix19_En18
  input [18:0] Wgt_7_415, // sfix19_En18
  input [18:0] Wgt_7_416, // sfix19_En18
  input [18:0] Wgt_7_417, // sfix19_En18
  input [18:0] Wgt_7_418, // sfix19_En18
  input [18:0] Wgt_7_419, // sfix19_En18
  input [18:0] Wgt_7_420, // sfix19_En18
  input [18:0] Wgt_7_421, // sfix19_En18
  input [18:0] Wgt_7_422, // sfix19_En18
  input [18:0] Wgt_7_423, // sfix19_En18
  input [18:0] Wgt_7_424, // sfix19_En18
  input [18:0] Wgt_7_425, // sfix19_En18
  input [18:0] Wgt_7_426, // sfix19_En18
  input [18:0] Wgt_7_427, // sfix19_En18
  input [18:0] Wgt_7_428, // sfix19_En18
  input [18:0] Wgt_7_429, // sfix19_En18
  input [18:0] Wgt_7_430, // sfix19_En18
  input [18:0] Wgt_7_431, // sfix19_En18
  input [18:0] Wgt_7_432, // sfix19_En18
  input [18:0] Wgt_7_433, // sfix19_En18
  input [18:0] Wgt_7_434, // sfix19_En18
  input [18:0] Wgt_7_435, // sfix19_En18
  input [18:0] Wgt_7_436, // sfix19_En18
  input [18:0] Wgt_7_437, // sfix19_En18
  input [18:0] Wgt_7_438, // sfix19_En18
  input [18:0] Wgt_7_439, // sfix19_En18
  input [18:0] Wgt_7_440, // sfix19_En18
  input [18:0] Wgt_7_441, // sfix19_En18
  input [18:0] Wgt_7_442, // sfix19_En18
  input [18:0] Wgt_7_443, // sfix19_En18
  input [18:0] Wgt_7_444, // sfix19_En18
  input [18:0] Wgt_7_445, // sfix19_En18
  input [18:0] Wgt_7_446, // sfix19_En18
  input [18:0] Wgt_7_447, // sfix19_En18
  input [18:0] Wgt_7_448, // sfix19_En18
  input [18:0] Wgt_7_449, // sfix19_En18
  input [18:0] Wgt_7_450, // sfix19_En18
  input [18:0] Wgt_7_451, // sfix19_En18
  input [18:0] Wgt_7_452, // sfix19_En18
  input [18:0] Wgt_7_453, // sfix19_En18
  input [18:0] Wgt_7_454, // sfix19_En18
  input [18:0] Wgt_7_455, // sfix19_En18
  input [18:0] Wgt_7_456, // sfix19_En18
  input [18:0] Wgt_7_457, // sfix19_En18
  input [18:0] Wgt_7_458, // sfix19_En18
  input [18:0] Wgt_7_459, // sfix19_En18
  input [18:0] Wgt_7_460, // sfix19_En18
  input [18:0] Wgt_7_461, // sfix19_En18
  input [18:0] Wgt_7_462, // sfix19_En18
  input [18:0] Wgt_7_463, // sfix19_En18
  input [18:0] Wgt_7_464, // sfix19_En18
  input [18:0] Wgt_7_465, // sfix19_En18
  input [18:0] Wgt_7_466, // sfix19_En18
  input [18:0] Wgt_7_467, // sfix19_En18
  input [18:0] Wgt_7_468, // sfix19_En18
  input [18:0] Wgt_7_469, // sfix19_En18
  input [18:0] Wgt_7_470, // sfix19_En18
  input [18:0] Wgt_7_471, // sfix19_En18
  input [18:0] Wgt_7_472, // sfix19_En18
  input [18:0] Wgt_7_473, // sfix19_En18
  input [18:0] Wgt_7_474, // sfix19_En18
  input [18:0] Wgt_7_475, // sfix19_En18
  input [18:0] Wgt_7_476, // sfix19_En18
  input [18:0] Wgt_7_477, // sfix19_En18
  input [18:0] Wgt_7_478, // sfix19_En18
  input [18:0] Wgt_7_479, // sfix19_En18
  input [18:0] Wgt_7_480, // sfix19_En18
  input [18:0] Wgt_7_481, // sfix19_En18
  input [18:0] Wgt_7_482, // sfix19_En18
  input [18:0] Wgt_7_483, // sfix19_En18
  input [18:0] Wgt_7_484, // sfix19_En18
  input [18:0] Wgt_7_485, // sfix19_En18
  input [18:0] Wgt_7_486, // sfix19_En18
  input [18:0] Wgt_7_487, // sfix19_En18
  input [18:0] Wgt_7_488, // sfix19_En18
  input [18:0] Wgt_7_489, // sfix19_En18
  input [18:0] Wgt_7_490, // sfix19_En18
  input [18:0] Wgt_7_491, // sfix19_En18
  input [18:0] Wgt_7_492, // sfix19_En18
  input [18:0] Wgt_7_493, // sfix19_En18
  input [18:0] Wgt_7_494, // sfix19_En18
  input [18:0] Wgt_7_495, // sfix19_En18
  input [18:0] Wgt_7_496, // sfix19_En18
  input [18:0] Wgt_7_497, // sfix19_En18
  input [18:0] Wgt_7_498, // sfix19_En18
  input [18:0] Wgt_7_499, // sfix19_En18
  input [18:0] Wgt_7_500, // sfix19_En18
  input [18:0] Wgt_7_501, // sfix19_En18
  input [18:0] Wgt_7_502, // sfix19_En18
  input [18:0] Wgt_7_503, // sfix19_En18
  input [18:0] Wgt_7_504, // sfix19_En18
  input [18:0] Wgt_7_505, // sfix19_En18
  input [18:0] Wgt_7_506, // sfix19_En18
  input [18:0] Wgt_7_507, // sfix19_En18
  input [18:0] Wgt_7_508, // sfix19_En18
  input [18:0] Wgt_7_509, // sfix19_En18
  input [18:0] Wgt_7_510, // sfix19_En18
  input [18:0] Wgt_7_511, // sfix19_En18
  input [18:0] Wgt_7_512, // sfix19_En18
  input [18:0] Wgt_7_513, // sfix19_En18
  input [18:0] Wgt_7_514, // sfix19_En18
  input [18:0] Wgt_7_515, // sfix19_En18
  input [18:0] Wgt_7_516, // sfix19_En18
  input [18:0] Wgt_7_517, // sfix19_En18
  input [18:0] Wgt_7_518, // sfix19_En18
  input [18:0] Wgt_7_519, // sfix19_En18
  input [18:0] Wgt_7_520, // sfix19_En18
  input [18:0] Wgt_7_521, // sfix19_En18
  input [18:0] Wgt_7_522, // sfix19_En18
  input [18:0] Wgt_7_523, // sfix19_En18
  input [18:0] Wgt_7_524, // sfix19_En18
  input [18:0] Wgt_7_525, // sfix19_En18
  input [18:0] Wgt_7_526, // sfix19_En18
  input [18:0] Wgt_7_527, // sfix19_En18
  input [18:0] Wgt_7_528, // sfix19_En18
  input [18:0] Wgt_7_529, // sfix19_En18
  input [18:0] Wgt_7_530, // sfix19_En18
  input [18:0] Wgt_7_531, // sfix19_En18
  input [18:0] Wgt_7_532, // sfix19_En18
  input [18:0] Wgt_7_533, // sfix19_En18
  input [18:0] Wgt_7_534, // sfix19_En18
  input [18:0] Wgt_7_535, // sfix19_En18
  input [18:0] Wgt_7_536, // sfix19_En18
  input [18:0] Wgt_7_537, // sfix19_En18
  input [18:0] Wgt_7_538, // sfix19_En18
  input [18:0] Wgt_7_539, // sfix19_En18
  input [18:0] Wgt_7_540, // sfix19_En18
  input [18:0] Wgt_7_541, // sfix19_En18
  input [18:0] Wgt_7_542, // sfix19_En18
  input [18:0] Wgt_7_543, // sfix19_En18
  input [18:0] Wgt_7_544, // sfix19_En18
  input [18:0] Wgt_7_545, // sfix19_En18
  input [18:0] Wgt_7_546, // sfix19_En18
  input [18:0] Wgt_7_547, // sfix19_En18
  input [18:0] Wgt_7_548, // sfix19_En18
  input [18:0] Wgt_7_549, // sfix19_En18
  input [18:0] Wgt_7_550, // sfix19_En18
  input [18:0] Wgt_7_551, // sfix19_En18
  input [18:0] Wgt_7_552, // sfix19_En18
  input [18:0] Wgt_7_553, // sfix19_En18
  input [18:0] Wgt_7_554, // sfix19_En18
  input [18:0] Wgt_7_555, // sfix19_En18
  input [18:0] Wgt_7_556, // sfix19_En18
  input [18:0] Wgt_7_557, // sfix19_En18
  input [18:0] Wgt_7_558, // sfix19_En18
  input [18:0] Wgt_7_559, // sfix19_En18
  input [18:0] Wgt_7_560, // sfix19_En18
  input [18:0] Wgt_7_561, // sfix19_En18
  input [18:0] Wgt_7_562, // sfix19_En18
  input [18:0] Wgt_7_563, // sfix19_En18
  input [18:0] Wgt_7_564, // sfix19_En18
  input [18:0] Wgt_7_565, // sfix19_En18
  input [18:0] Wgt_7_566, // sfix19_En18
  input [18:0] Wgt_7_567, // sfix19_En18
  input [18:0] Wgt_7_568, // sfix19_En18
  input [18:0] Wgt_7_569, // sfix19_En18
  input [18:0] Wgt_7_570, // sfix19_En18
  input [18:0] Wgt_7_571, // sfix19_En18
  input [18:0] Wgt_7_572, // sfix19_En18
  input [18:0] Wgt_7_573, // sfix19_En18
  input [18:0] Wgt_7_574, // sfix19_En18
  input [18:0] Wgt_7_575, // sfix19_En18
  input [18:0] Wgt_7_576, // sfix19_En18
  input [18:0] Wgt_7_577, // sfix19_En18
  input [18:0] Wgt_7_578, // sfix19_En18
  input [18:0] Wgt_7_579, // sfix19_En18
  input [18:0] Wgt_7_580, // sfix19_En18
  input [18:0] Wgt_7_581, // sfix19_En18
  input [18:0] Wgt_7_582, // sfix19_En18
  input [18:0] Wgt_7_583, // sfix19_En18
  input [18:0] Wgt_7_584, // sfix19_En18
  input [18:0] Wgt_7_585, // sfix19_En18
  input [18:0] Wgt_7_586, // sfix19_En18
  input [18:0] Wgt_7_587, // sfix19_En18
  input [18:0] Wgt_7_588, // sfix19_En18
  input [18:0] Wgt_7_589, // sfix19_En18
  input [18:0] Wgt_7_590, // sfix19_En18
  input [18:0] Wgt_7_591, // sfix19_En18
  input [18:0] Wgt_7_592, // sfix19_En18
  input [18:0] Wgt_7_593, // sfix19_En18
  input [18:0] Wgt_7_594, // sfix19_En18
  input [18:0] Wgt_7_595, // sfix19_En18
  input [18:0] Wgt_7_596, // sfix19_En18
  input [18:0] Wgt_7_597, // sfix19_En18
  input [18:0] Wgt_7_598, // sfix19_En18
  input [18:0] Wgt_7_599, // sfix19_En18
  input [18:0] Wgt_7_600, // sfix19_En18
  input [18:0] Wgt_7_601, // sfix19_En18
  input [18:0] Wgt_7_602, // sfix19_En18
  input [18:0] Wgt_7_603, // sfix19_En18
  input [18:0] Wgt_7_604, // sfix19_En18
  input [18:0] Wgt_7_605, // sfix19_En18
  input [18:0] Wgt_7_606, // sfix19_En18
  input [18:0] Wgt_7_607, // sfix19_En18
  input [18:0] Wgt_7_608, // sfix19_En18
  input [18:0] Wgt_7_609, // sfix19_En18
  input [18:0] Wgt_7_610, // sfix19_En18
  input [18:0] Wgt_7_611, // sfix19_En18
  input [18:0] Wgt_7_612, // sfix19_En18
  input [18:0] Wgt_7_613, // sfix19_En18
  input [18:0] Wgt_7_614, // sfix19_En18
  input [18:0] Wgt_7_615, // sfix19_En18
  input [18:0] Wgt_7_616, // sfix19_En18
  input [18:0] Wgt_7_617, // sfix19_En18
  input [18:0] Wgt_7_618, // sfix19_En18
  input [18:0] Wgt_7_619, // sfix19_En18
  input [18:0] Wgt_7_620, // sfix19_En18
  input [18:0] Wgt_7_621, // sfix19_En18
  input [18:0] Wgt_7_622, // sfix19_En18
  input [18:0] Wgt_7_623, // sfix19_En18
  input [18:0] Wgt_7_624, // sfix19_En18
  input [18:0] Wgt_7_625, // sfix19_En18
  input [18:0] Wgt_7_626, // sfix19_En18
  input [18:0] Wgt_7_627, // sfix19_En18
  input [18:0] Wgt_7_628, // sfix19_En18
  input [18:0] Wgt_7_629, // sfix19_En18
  input [18:0] Wgt_7_630, // sfix19_En18
  input [18:0] Wgt_7_631, // sfix19_En18
  input [18:0] Wgt_7_632, // sfix19_En18
  input [18:0] Wgt_7_633, // sfix19_En18
  input [18:0] Wgt_7_634, // sfix19_En18
  input [18:0] Wgt_7_635, // sfix19_En18
  input [18:0] Wgt_7_636, // sfix19_En18
  input [18:0] Wgt_7_637, // sfix19_En18
  input [18:0] Wgt_7_638, // sfix19_En18
  input [18:0] Wgt_7_639, // sfix19_En18
  input [18:0] Wgt_7_640, // sfix19_En18
  input [18:0] Wgt_7_641, // sfix19_En18
  input [18:0] Wgt_7_642, // sfix19_En18
  input [18:0] Wgt_7_643, // sfix19_En18
  input [18:0] Wgt_7_644, // sfix19_En18
  input [18:0] Wgt_7_645, // sfix19_En18
  input [18:0] Wgt_7_646, // sfix19_En18
  input [18:0] Wgt_7_647, // sfix19_En18
  input [18:0] Wgt_7_648, // sfix19_En18
  input [18:0] Wgt_7_649, // sfix19_En18
  input [18:0] Wgt_7_650, // sfix19_En18
  input [18:0] Wgt_7_651, // sfix19_En18
  input [18:0] Wgt_7_652, // sfix19_En18
  input [18:0] Wgt_7_653, // sfix19_En18
  input [18:0] Wgt_7_654, // sfix19_En18
  input [18:0] Wgt_7_655, // sfix19_En18
  input [18:0] Wgt_7_656, // sfix19_En18
  input [18:0] Wgt_7_657, // sfix19_En18
  input [18:0] Wgt_7_658, // sfix19_En18
  input [18:0] Wgt_7_659, // sfix19_En18
  input [18:0] Wgt_7_660, // sfix19_En18
  input [18:0] Wgt_7_661, // sfix19_En18
  input [18:0] Wgt_7_662, // sfix19_En18
  input [18:0] Wgt_7_663, // sfix19_En18
  input [18:0] Wgt_7_664, // sfix19_En18
  input [18:0] Wgt_7_665, // sfix19_En18
  input [18:0] Wgt_7_666, // sfix19_En18
  input [18:0] Wgt_7_667, // sfix19_En18
  input [18:0] Wgt_7_668, // sfix19_En18
  input [18:0] Wgt_7_669, // sfix19_En18
  input [18:0] Wgt_7_670, // sfix19_En18
  input [18:0] Wgt_7_671, // sfix19_En18
  input [18:0] Wgt_7_672, // sfix19_En18
  input [18:0] Wgt_7_673, // sfix19_En18
  input [18:0] Wgt_7_674, // sfix19_En18
  input [18:0] Wgt_7_675, // sfix19_En18
  input [18:0] Wgt_7_676, // sfix19_En18
  input [18:0] Wgt_7_677, // sfix19_En18
  input [18:0] Wgt_7_678, // sfix19_En18
  input [18:0] Wgt_7_679, // sfix19_En18
  input [18:0] Wgt_7_680, // sfix19_En18
  input [18:0] Wgt_7_681, // sfix19_En18
  input [18:0] Wgt_7_682, // sfix19_En18
  input [18:0] Wgt_7_683, // sfix19_En18
  input [18:0] Wgt_7_684, // sfix19_En18
  input [18:0] Wgt_7_685, // sfix19_En18
  input [18:0] Wgt_7_686, // sfix19_En18
  input [18:0] Wgt_7_687, // sfix19_En18
  input [18:0] Wgt_7_688, // sfix19_En18
  input [18:0] Wgt_7_689, // sfix19_En18
  input [18:0] Wgt_7_690, // sfix19_En18
  input [18:0] Wgt_7_691, // sfix19_En18
  input [18:0] Wgt_7_692, // sfix19_En18
  input [18:0] Wgt_7_693, // sfix19_En18
  input [18:0] Wgt_7_694, // sfix19_En18
  input [18:0] Wgt_7_695, // sfix19_En18
  input [18:0] Wgt_7_696, // sfix19_En18
  input [18:0] Wgt_7_697, // sfix19_En18
  input [18:0] Wgt_7_698, // sfix19_En18
  input [18:0] Wgt_7_699, // sfix19_En18
  input [18:0] Wgt_7_700, // sfix19_En18
  input [18:0] Wgt_7_701, // sfix19_En18
  input [18:0] Wgt_7_702, // sfix19_En18
  input [18:0] Wgt_7_703, // sfix19_En18
  input [18:0] Wgt_7_704, // sfix19_En18
  input [18:0] Wgt_7_705, // sfix19_En18
  input [18:0] Wgt_7_706, // sfix19_En18
  input [18:0] Wgt_7_707, // sfix19_En18
  input [18:0] Wgt_7_708, // sfix19_En18
  input [18:0] Wgt_7_709, // sfix19_En18
  input [18:0] Wgt_7_710, // sfix19_En18
  input [18:0] Wgt_7_711, // sfix19_En18
  input [18:0] Wgt_7_712, // sfix19_En18
  input [18:0] Wgt_7_713, // sfix19_En18
  input [18:0] Wgt_7_714, // sfix19_En18
  input [18:0] Wgt_7_715, // sfix19_En18
  input [18:0] Wgt_7_716, // sfix19_En18
  input [18:0] Wgt_7_717, // sfix19_En18
  input [18:0] Wgt_7_718, // sfix19_En18
  input [18:0] Wgt_7_719, // sfix19_En18
  input [18:0] Wgt_7_720, // sfix19_En18
  input [18:0] Wgt_7_721, // sfix19_En18
  input [18:0] Wgt_7_722, // sfix19_En18
  input [18:0] Wgt_7_723, // sfix19_En18
  input [18:0] Wgt_7_724, // sfix19_En18
  input [18:0] Wgt_7_725, // sfix19_En18
  input [18:0] Wgt_7_726, // sfix19_En18
  input [18:0] Wgt_7_727, // sfix19_En18
  input [18:0] Wgt_7_728, // sfix19_En18
  input [18:0] Wgt_7_729, // sfix19_En18
  input [18:0] Wgt_7_730, // sfix19_En18
  input [18:0] Wgt_7_731, // sfix19_En18
  input [18:0] Wgt_7_732, // sfix19_En18
  input [18:0] Wgt_7_733, // sfix19_En18
  input [18:0] Wgt_7_734, // sfix19_En18
  input [18:0] Wgt_7_735, // sfix19_En18
  input [18:0] Wgt_7_736, // sfix19_En18
  input [18:0] Wgt_7_737, // sfix19_En18
  input [18:0] Wgt_7_738, // sfix19_En18
  input [18:0] Wgt_7_739, // sfix19_En18
  input [18:0] Wgt_7_740, // sfix19_En18
  input [18:0] Wgt_7_741, // sfix19_En18
  input [18:0] Wgt_7_742, // sfix19_En18
  input [18:0] Wgt_7_743, // sfix19_En18
  input [18:0] Wgt_7_744, // sfix19_En18
  input [18:0] Wgt_7_745, // sfix19_En18
  input [18:0] Wgt_7_746, // sfix19_En18
  input [18:0] Wgt_7_747, // sfix19_En18
  input [18:0] Wgt_7_748, // sfix19_En18
  input [18:0] Wgt_7_749, // sfix19_En18
  input [18:0] Wgt_7_750, // sfix19_En18
  input [18:0] Wgt_7_751, // sfix19_En18
  input [18:0] Wgt_7_752, // sfix19_En18
  input [18:0] Wgt_7_753, // sfix19_En18
  input [18:0] Wgt_7_754, // sfix19_En18
  input [18:0] Wgt_7_755, // sfix19_En18
  input [18:0] Wgt_7_756, // sfix19_En18
  input [18:0] Wgt_7_757, // sfix19_En18
  input [18:0] Wgt_7_758, // sfix19_En18
  input [18:0] Wgt_7_759, // sfix19_En18
  input [18:0] Wgt_7_760, // sfix19_En18
  input [18:0] Wgt_7_761, // sfix19_En18
  input [18:0] Wgt_7_762, // sfix19_En18
  input [18:0] Wgt_7_763, // sfix19_En18
  input [18:0] Wgt_7_764, // sfix19_En18
  input [18:0] Wgt_7_765, // sfix19_En18
  input [18:0] Wgt_7_766, // sfix19_En18
  input [18:0] Wgt_7_767, // sfix19_En18
  input [18:0] Wgt_7_768, // sfix19_En18
  input [18:0] Wgt_7_769, // sfix19_En18
  input [18:0] Wgt_7_770, // sfix19_En18
  input [18:0] Wgt_7_771, // sfix19_En18
  input [18:0] Wgt_7_772, // sfix19_En18
  input [18:0] Wgt_7_773, // sfix19_En18
  input [18:0] Wgt_7_774, // sfix19_En18
  input [18:0] Wgt_7_775, // sfix19_En18
  input [18:0] Wgt_7_776, // sfix19_En18
  input [18:0] Wgt_7_777, // sfix19_En18
  input [18:0] Wgt_7_778, // sfix19_En18
  input [18:0] Wgt_7_779, // sfix19_En18
  input [18:0] Wgt_7_780, // sfix19_En18
  input [18:0] Wgt_7_781, // sfix19_En18
  input [18:0] Wgt_7_782, // sfix19_En18
  input [18:0] Wgt_7_783, // sfix19_En18
  input [18:0] Wgt_7_784, // sfix19_En18
  input [18:0] Wgt_8_0, // sfix19_En18
  input [18:0] Wgt_8_1, // sfix19_En18
  input [18:0] Wgt_8_2, // sfix19_En18
  input [18:0] Wgt_8_3, // sfix19_En18
  input [18:0] Wgt_8_4, // sfix19_En18
  input [18:0] Wgt_8_5, // sfix19_En18
  input [18:0] Wgt_8_6, // sfix19_En18
  input [18:0] Wgt_8_7, // sfix19_En18
  input [18:0] Wgt_8_8, // sfix19_En18
  input [18:0] Wgt_8_9, // sfix19_En18
  input [18:0] Wgt_8_10, // sfix19_En18
  input [18:0] Wgt_8_11, // sfix19_En18
  input [18:0] Wgt_8_12, // sfix19_En18
  input [18:0] Wgt_8_13, // sfix19_En18
  input [18:0] Wgt_8_14, // sfix19_En18
  input [18:0] Wgt_8_15, // sfix19_En18
  input [18:0] Wgt_8_16, // sfix19_En18
  input [18:0] Wgt_8_17, // sfix19_En18
  input [18:0] Wgt_8_18, // sfix19_En18
  input [18:0] Wgt_8_19, // sfix19_En18
  input [18:0] Wgt_8_20, // sfix19_En18
  input [18:0] Wgt_8_21, // sfix19_En18
  input [18:0] Wgt_8_22, // sfix19_En18
  input [18:0] Wgt_8_23, // sfix19_En18
  input [18:0] Wgt_8_24, // sfix19_En18
  input [18:0] Wgt_8_25, // sfix19_En18
  input [18:0] Wgt_8_26, // sfix19_En18
  input [18:0] Wgt_8_27, // sfix19_En18
  input [18:0] Wgt_8_28, // sfix19_En18
  input [18:0] Wgt_8_29, // sfix19_En18
  input [18:0] Wgt_8_30, // sfix19_En18
  input [18:0] Wgt_8_31, // sfix19_En18
  input [18:0] Wgt_8_32, // sfix19_En18
  input [18:0] Wgt_8_33, // sfix19_En18
  input [18:0] Wgt_8_34, // sfix19_En18
  input [18:0] Wgt_8_35, // sfix19_En18
  input [18:0] Wgt_8_36, // sfix19_En18
  input [18:0] Wgt_8_37, // sfix19_En18
  input [18:0] Wgt_8_38, // sfix19_En18
  input [18:0] Wgt_8_39, // sfix19_En18
  input [18:0] Wgt_8_40, // sfix19_En18
  input [18:0] Wgt_8_41, // sfix19_En18
  input [18:0] Wgt_8_42, // sfix19_En18
  input [18:0] Wgt_8_43, // sfix19_En18
  input [18:0] Wgt_8_44, // sfix19_En18
  input [18:0] Wgt_8_45, // sfix19_En18
  input [18:0] Wgt_8_46, // sfix19_En18
  input [18:0] Wgt_8_47, // sfix19_En18
  input [18:0] Wgt_8_48, // sfix19_En18
  input [18:0] Wgt_8_49, // sfix19_En18
  input [18:0] Wgt_8_50, // sfix19_En18
  input [18:0] Wgt_8_51, // sfix19_En18
  input [18:0] Wgt_8_52, // sfix19_En18
  input [18:0] Wgt_8_53, // sfix19_En18
  input [18:0] Wgt_8_54, // sfix19_En18
  input [18:0] Wgt_8_55, // sfix19_En18
  input [18:0] Wgt_8_56, // sfix19_En18
  input [18:0] Wgt_8_57, // sfix19_En18
  input [18:0] Wgt_8_58, // sfix19_En18
  input [18:0] Wgt_8_59, // sfix19_En18
  input [18:0] Wgt_8_60, // sfix19_En18
  input [18:0] Wgt_8_61, // sfix19_En18
  input [18:0] Wgt_8_62, // sfix19_En18
  input [18:0] Wgt_8_63, // sfix19_En18
  input [18:0] Wgt_8_64, // sfix19_En18
  input [18:0] Wgt_8_65, // sfix19_En18
  input [18:0] Wgt_8_66, // sfix19_En18
  input [18:0] Wgt_8_67, // sfix19_En18
  input [18:0] Wgt_8_68, // sfix19_En18
  input [18:0] Wgt_8_69, // sfix19_En18
  input [18:0] Wgt_8_70, // sfix19_En18
  input [18:0] Wgt_8_71, // sfix19_En18
  input [18:0] Wgt_8_72, // sfix19_En18
  input [18:0] Wgt_8_73, // sfix19_En18
  input [18:0] Wgt_8_74, // sfix19_En18
  input [18:0] Wgt_8_75, // sfix19_En18
  input [18:0] Wgt_8_76, // sfix19_En18
  input [18:0] Wgt_8_77, // sfix19_En18
  input [18:0] Wgt_8_78, // sfix19_En18
  input [18:0] Wgt_8_79, // sfix19_En18
  input [18:0] Wgt_8_80, // sfix19_En18
  input [18:0] Wgt_8_81, // sfix19_En18
  input [18:0] Wgt_8_82, // sfix19_En18
  input [18:0] Wgt_8_83, // sfix19_En18
  input [18:0] Wgt_8_84, // sfix19_En18
  input [18:0] Wgt_8_85, // sfix19_En18
  input [18:0] Wgt_8_86, // sfix19_En18
  input [18:0] Wgt_8_87, // sfix19_En18
  input [18:0] Wgt_8_88, // sfix19_En18
  input [18:0] Wgt_8_89, // sfix19_En18
  input [18:0] Wgt_8_90, // sfix19_En18
  input [18:0] Wgt_8_91, // sfix19_En18
  input [18:0] Wgt_8_92, // sfix19_En18
  input [18:0] Wgt_8_93, // sfix19_En18
  input [18:0] Wgt_8_94, // sfix19_En18
  input [18:0] Wgt_8_95, // sfix19_En18
  input [18:0] Wgt_8_96, // sfix19_En18
  input [18:0] Wgt_8_97, // sfix19_En18
  input [18:0] Wgt_8_98, // sfix19_En18
  input [18:0] Wgt_8_99, // sfix19_En18
  input [18:0] Wgt_8_100, // sfix19_En18
  input [18:0] Wgt_8_101, // sfix19_En18
  input [18:0] Wgt_8_102, // sfix19_En18
  input [18:0] Wgt_8_103, // sfix19_En18
  input [18:0] Wgt_8_104, // sfix19_En18
  input [18:0] Wgt_8_105, // sfix19_En18
  input [18:0] Wgt_8_106, // sfix19_En18
  input [18:0] Wgt_8_107, // sfix19_En18
  input [18:0] Wgt_8_108, // sfix19_En18
  input [18:0] Wgt_8_109, // sfix19_En18
  input [18:0] Wgt_8_110, // sfix19_En18
  input [18:0] Wgt_8_111, // sfix19_En18
  input [18:0] Wgt_8_112, // sfix19_En18
  input [18:0] Wgt_8_113, // sfix19_En18
  input [18:0] Wgt_8_114, // sfix19_En18
  input [18:0] Wgt_8_115, // sfix19_En18
  input [18:0] Wgt_8_116, // sfix19_En18
  input [18:0] Wgt_8_117, // sfix19_En18
  input [18:0] Wgt_8_118, // sfix19_En18
  input [18:0] Wgt_8_119, // sfix19_En18
  input [18:0] Wgt_8_120, // sfix19_En18
  input [18:0] Wgt_8_121, // sfix19_En18
  input [18:0] Wgt_8_122, // sfix19_En18
  input [18:0] Wgt_8_123, // sfix19_En18
  input [18:0] Wgt_8_124, // sfix19_En18
  input [18:0] Wgt_8_125, // sfix19_En18
  input [18:0] Wgt_8_126, // sfix19_En18
  input [18:0] Wgt_8_127, // sfix19_En18
  input [18:0] Wgt_8_128, // sfix19_En18
  input [18:0] Wgt_8_129, // sfix19_En18
  input [18:0] Wgt_8_130, // sfix19_En18
  input [18:0] Wgt_8_131, // sfix19_En18
  input [18:0] Wgt_8_132, // sfix19_En18
  input [18:0] Wgt_8_133, // sfix19_En18
  input [18:0] Wgt_8_134, // sfix19_En18
  input [18:0] Wgt_8_135, // sfix19_En18
  input [18:0] Wgt_8_136, // sfix19_En18
  input [18:0] Wgt_8_137, // sfix19_En18
  input [18:0] Wgt_8_138, // sfix19_En18
  input [18:0] Wgt_8_139, // sfix19_En18
  input [18:0] Wgt_8_140, // sfix19_En18
  input [18:0] Wgt_8_141, // sfix19_En18
  input [18:0] Wgt_8_142, // sfix19_En18
  input [18:0] Wgt_8_143, // sfix19_En18
  input [18:0] Wgt_8_144, // sfix19_En18
  input [18:0] Wgt_8_145, // sfix19_En18
  input [18:0] Wgt_8_146, // sfix19_En18
  input [18:0] Wgt_8_147, // sfix19_En18
  input [18:0] Wgt_8_148, // sfix19_En18
  input [18:0] Wgt_8_149, // sfix19_En18
  input [18:0] Wgt_8_150, // sfix19_En18
  input [18:0] Wgt_8_151, // sfix19_En18
  input [18:0] Wgt_8_152, // sfix19_En18
  input [18:0] Wgt_8_153, // sfix19_En18
  input [18:0] Wgt_8_154, // sfix19_En18
  input [18:0] Wgt_8_155, // sfix19_En18
  input [18:0] Wgt_8_156, // sfix19_En18
  input [18:0] Wgt_8_157, // sfix19_En18
  input [18:0] Wgt_8_158, // sfix19_En18
  input [18:0] Wgt_8_159, // sfix19_En18
  input [18:0] Wgt_8_160, // sfix19_En18
  input [18:0] Wgt_8_161, // sfix19_En18
  input [18:0] Wgt_8_162, // sfix19_En18
  input [18:0] Wgt_8_163, // sfix19_En18
  input [18:0] Wgt_8_164, // sfix19_En18
  input [18:0] Wgt_8_165, // sfix19_En18
  input [18:0] Wgt_8_166, // sfix19_En18
  input [18:0] Wgt_8_167, // sfix19_En18
  input [18:0] Wgt_8_168, // sfix19_En18
  input [18:0] Wgt_8_169, // sfix19_En18
  input [18:0] Wgt_8_170, // sfix19_En18
  input [18:0] Wgt_8_171, // sfix19_En18
  input [18:0] Wgt_8_172, // sfix19_En18
  input [18:0] Wgt_8_173, // sfix19_En18
  input [18:0] Wgt_8_174, // sfix19_En18
  input [18:0] Wgt_8_175, // sfix19_En18
  input [18:0] Wgt_8_176, // sfix19_En18
  input [18:0] Wgt_8_177, // sfix19_En18
  input [18:0] Wgt_8_178, // sfix19_En18
  input [18:0] Wgt_8_179, // sfix19_En18
  input [18:0] Wgt_8_180, // sfix19_En18
  input [18:0] Wgt_8_181, // sfix19_En18
  input [18:0] Wgt_8_182, // sfix19_En18
  input [18:0] Wgt_8_183, // sfix19_En18
  input [18:0] Wgt_8_184, // sfix19_En18
  input [18:0] Wgt_8_185, // sfix19_En18
  input [18:0] Wgt_8_186, // sfix19_En18
  input [18:0] Wgt_8_187, // sfix19_En18
  input [18:0] Wgt_8_188, // sfix19_En18
  input [18:0] Wgt_8_189, // sfix19_En18
  input [18:0] Wgt_8_190, // sfix19_En18
  input [18:0] Wgt_8_191, // sfix19_En18
  input [18:0] Wgt_8_192, // sfix19_En18
  input [18:0] Wgt_8_193, // sfix19_En18
  input [18:0] Wgt_8_194, // sfix19_En18
  input [18:0] Wgt_8_195, // sfix19_En18
  input [18:0] Wgt_8_196, // sfix19_En18
  input [18:0] Wgt_8_197, // sfix19_En18
  input [18:0] Wgt_8_198, // sfix19_En18
  input [18:0] Wgt_8_199, // sfix19_En18
  input [18:0] Wgt_8_200, // sfix19_En18
  input [18:0] Wgt_8_201, // sfix19_En18
  input [18:0] Wgt_8_202, // sfix19_En18
  input [18:0] Wgt_8_203, // sfix19_En18
  input [18:0] Wgt_8_204, // sfix19_En18
  input [18:0] Wgt_8_205, // sfix19_En18
  input [18:0] Wgt_8_206, // sfix19_En18
  input [18:0] Wgt_8_207, // sfix19_En18
  input [18:0] Wgt_8_208, // sfix19_En18
  input [18:0] Wgt_8_209, // sfix19_En18
  input [18:0] Wgt_8_210, // sfix19_En18
  input [18:0] Wgt_8_211, // sfix19_En18
  input [18:0] Wgt_8_212, // sfix19_En18
  input [18:0] Wgt_8_213, // sfix19_En18
  input [18:0] Wgt_8_214, // sfix19_En18
  input [18:0] Wgt_8_215, // sfix19_En18
  input [18:0] Wgt_8_216, // sfix19_En18
  input [18:0] Wgt_8_217, // sfix19_En18
  input [18:0] Wgt_8_218, // sfix19_En18
  input [18:0] Wgt_8_219, // sfix19_En18
  input [18:0] Wgt_8_220, // sfix19_En18
  input [18:0] Wgt_8_221, // sfix19_En18
  input [18:0] Wgt_8_222, // sfix19_En18
  input [18:0] Wgt_8_223, // sfix19_En18
  input [18:0] Wgt_8_224, // sfix19_En18
  input [18:0] Wgt_8_225, // sfix19_En18
  input [18:0] Wgt_8_226, // sfix19_En18
  input [18:0] Wgt_8_227, // sfix19_En18
  input [18:0] Wgt_8_228, // sfix19_En18
  input [18:0] Wgt_8_229, // sfix19_En18
  input [18:0] Wgt_8_230, // sfix19_En18
  input [18:0] Wgt_8_231, // sfix19_En18
  input [18:0] Wgt_8_232, // sfix19_En18
  input [18:0] Wgt_8_233, // sfix19_En18
  input [18:0] Wgt_8_234, // sfix19_En18
  input [18:0] Wgt_8_235, // sfix19_En18
  input [18:0] Wgt_8_236, // sfix19_En18
  input [18:0] Wgt_8_237, // sfix19_En18
  input [18:0] Wgt_8_238, // sfix19_En18
  input [18:0] Wgt_8_239, // sfix19_En18
  input [18:0] Wgt_8_240, // sfix19_En18
  input [18:0] Wgt_8_241, // sfix19_En18
  input [18:0] Wgt_8_242, // sfix19_En18
  input [18:0] Wgt_8_243, // sfix19_En18
  input [18:0] Wgt_8_244, // sfix19_En18
  input [18:0] Wgt_8_245, // sfix19_En18
  input [18:0] Wgt_8_246, // sfix19_En18
  input [18:0] Wgt_8_247, // sfix19_En18
  input [18:0] Wgt_8_248, // sfix19_En18
  input [18:0] Wgt_8_249, // sfix19_En18
  input [18:0] Wgt_8_250, // sfix19_En18
  input [18:0] Wgt_8_251, // sfix19_En18
  input [18:0] Wgt_8_252, // sfix19_En18
  input [18:0] Wgt_8_253, // sfix19_En18
  input [18:0] Wgt_8_254, // sfix19_En18
  input [18:0] Wgt_8_255, // sfix19_En18
  input [18:0] Wgt_8_256, // sfix19_En18
  input [18:0] Wgt_8_257, // sfix19_En18
  input [18:0] Wgt_8_258, // sfix19_En18
  input [18:0] Wgt_8_259, // sfix19_En18
  input [18:0] Wgt_8_260, // sfix19_En18
  input [18:0] Wgt_8_261, // sfix19_En18
  input [18:0] Wgt_8_262, // sfix19_En18
  input [18:0] Wgt_8_263, // sfix19_En18
  input [18:0] Wgt_8_264, // sfix19_En18
  input [18:0] Wgt_8_265, // sfix19_En18
  input [18:0] Wgt_8_266, // sfix19_En18
  input [18:0] Wgt_8_267, // sfix19_En18
  input [18:0] Wgt_8_268, // sfix19_En18
  input [18:0] Wgt_8_269, // sfix19_En18
  input [18:0] Wgt_8_270, // sfix19_En18
  input [18:0] Wgt_8_271, // sfix19_En18
  input [18:0] Wgt_8_272, // sfix19_En18
  input [18:0] Wgt_8_273, // sfix19_En18
  input [18:0] Wgt_8_274, // sfix19_En18
  input [18:0] Wgt_8_275, // sfix19_En18
  input [18:0] Wgt_8_276, // sfix19_En18
  input [18:0] Wgt_8_277, // sfix19_En18
  input [18:0] Wgt_8_278, // sfix19_En18
  input [18:0] Wgt_8_279, // sfix19_En18
  input [18:0] Wgt_8_280, // sfix19_En18
  input [18:0] Wgt_8_281, // sfix19_En18
  input [18:0] Wgt_8_282, // sfix19_En18
  input [18:0] Wgt_8_283, // sfix19_En18
  input [18:0] Wgt_8_284, // sfix19_En18
  input [18:0] Wgt_8_285, // sfix19_En18
  input [18:0] Wgt_8_286, // sfix19_En18
  input [18:0] Wgt_8_287, // sfix19_En18
  input [18:0] Wgt_8_288, // sfix19_En18
  input [18:0] Wgt_8_289, // sfix19_En18
  input [18:0] Wgt_8_290, // sfix19_En18
  input [18:0] Wgt_8_291, // sfix19_En18
  input [18:0] Wgt_8_292, // sfix19_En18
  input [18:0] Wgt_8_293, // sfix19_En18
  input [18:0] Wgt_8_294, // sfix19_En18
  input [18:0] Wgt_8_295, // sfix19_En18
  input [18:0] Wgt_8_296, // sfix19_En18
  input [18:0] Wgt_8_297, // sfix19_En18
  input [18:0] Wgt_8_298, // sfix19_En18
  input [18:0] Wgt_8_299, // sfix19_En18
  input [18:0] Wgt_8_300, // sfix19_En18
  input [18:0] Wgt_8_301, // sfix19_En18
  input [18:0] Wgt_8_302, // sfix19_En18
  input [18:0] Wgt_8_303, // sfix19_En18
  input [18:0] Wgt_8_304, // sfix19_En18
  input [18:0] Wgt_8_305, // sfix19_En18
  input [18:0] Wgt_8_306, // sfix19_En18
  input [18:0] Wgt_8_307, // sfix19_En18
  input [18:0] Wgt_8_308, // sfix19_En18
  input [18:0] Wgt_8_309, // sfix19_En18
  input [18:0] Wgt_8_310, // sfix19_En18
  input [18:0] Wgt_8_311, // sfix19_En18
  input [18:0] Wgt_8_312, // sfix19_En18
  input [18:0] Wgt_8_313, // sfix19_En18
  input [18:0] Wgt_8_314, // sfix19_En18
  input [18:0] Wgt_8_315, // sfix19_En18
  input [18:0] Wgt_8_316, // sfix19_En18
  input [18:0] Wgt_8_317, // sfix19_En18
  input [18:0] Wgt_8_318, // sfix19_En18
  input [18:0] Wgt_8_319, // sfix19_En18
  input [18:0] Wgt_8_320, // sfix19_En18
  input [18:0] Wgt_8_321, // sfix19_En18
  input [18:0] Wgt_8_322, // sfix19_En18
  input [18:0] Wgt_8_323, // sfix19_En18
  input [18:0] Wgt_8_324, // sfix19_En18
  input [18:0] Wgt_8_325, // sfix19_En18
  input [18:0] Wgt_8_326, // sfix19_En18
  input [18:0] Wgt_8_327, // sfix19_En18
  input [18:0] Wgt_8_328, // sfix19_En18
  input [18:0] Wgt_8_329, // sfix19_En18
  input [18:0] Wgt_8_330, // sfix19_En18
  input [18:0] Wgt_8_331, // sfix19_En18
  input [18:0] Wgt_8_332, // sfix19_En18
  input [18:0] Wgt_8_333, // sfix19_En18
  input [18:0] Wgt_8_334, // sfix19_En18
  input [18:0] Wgt_8_335, // sfix19_En18
  input [18:0] Wgt_8_336, // sfix19_En18
  input [18:0] Wgt_8_337, // sfix19_En18
  input [18:0] Wgt_8_338, // sfix19_En18
  input [18:0] Wgt_8_339, // sfix19_En18
  input [18:0] Wgt_8_340, // sfix19_En18
  input [18:0] Wgt_8_341, // sfix19_En18
  input [18:0] Wgt_8_342, // sfix19_En18
  input [18:0] Wgt_8_343, // sfix19_En18
  input [18:0] Wgt_8_344, // sfix19_En18
  input [18:0] Wgt_8_345, // sfix19_En18
  input [18:0] Wgt_8_346, // sfix19_En18
  input [18:0] Wgt_8_347, // sfix19_En18
  input [18:0] Wgt_8_348, // sfix19_En18
  input [18:0] Wgt_8_349, // sfix19_En18
  input [18:0] Wgt_8_350, // sfix19_En18
  input [18:0] Wgt_8_351, // sfix19_En18
  input [18:0] Wgt_8_352, // sfix19_En18
  input [18:0] Wgt_8_353, // sfix19_En18
  input [18:0] Wgt_8_354, // sfix19_En18
  input [18:0] Wgt_8_355, // sfix19_En18
  input [18:0] Wgt_8_356, // sfix19_En18
  input [18:0] Wgt_8_357, // sfix19_En18
  input [18:0] Wgt_8_358, // sfix19_En18
  input [18:0] Wgt_8_359, // sfix19_En18
  input [18:0] Wgt_8_360, // sfix19_En18
  input [18:0] Wgt_8_361, // sfix19_En18
  input [18:0] Wgt_8_362, // sfix19_En18
  input [18:0] Wgt_8_363, // sfix19_En18
  input [18:0] Wgt_8_364, // sfix19_En18
  input [18:0] Wgt_8_365, // sfix19_En18
  input [18:0] Wgt_8_366, // sfix19_En18
  input [18:0] Wgt_8_367, // sfix19_En18
  input [18:0] Wgt_8_368, // sfix19_En18
  input [18:0] Wgt_8_369, // sfix19_En18
  input [18:0] Wgt_8_370, // sfix19_En18
  input [18:0] Wgt_8_371, // sfix19_En18
  input [18:0] Wgt_8_372, // sfix19_En18
  input [18:0] Wgt_8_373, // sfix19_En18
  input [18:0] Wgt_8_374, // sfix19_En18
  input [18:0] Wgt_8_375, // sfix19_En18
  input [18:0] Wgt_8_376, // sfix19_En18
  input [18:0] Wgt_8_377, // sfix19_En18
  input [18:0] Wgt_8_378, // sfix19_En18
  input [18:0] Wgt_8_379, // sfix19_En18
  input [18:0] Wgt_8_380, // sfix19_En18
  input [18:0] Wgt_8_381, // sfix19_En18
  input [18:0] Wgt_8_382, // sfix19_En18
  input [18:0] Wgt_8_383, // sfix19_En18
  input [18:0] Wgt_8_384, // sfix19_En18
  input [18:0] Wgt_8_385, // sfix19_En18
  input [18:0] Wgt_8_386, // sfix19_En18
  input [18:0] Wgt_8_387, // sfix19_En18
  input [18:0] Wgt_8_388, // sfix19_En18
  input [18:0] Wgt_8_389, // sfix19_En18
  input [18:0] Wgt_8_390, // sfix19_En18
  input [18:0] Wgt_8_391, // sfix19_En18
  input [18:0] Wgt_8_392, // sfix19_En18
  input [18:0] Wgt_8_393, // sfix19_En18
  input [18:0] Wgt_8_394, // sfix19_En18
  input [18:0] Wgt_8_395, // sfix19_En18
  input [18:0] Wgt_8_396, // sfix19_En18
  input [18:0] Wgt_8_397, // sfix19_En18
  input [18:0] Wgt_8_398, // sfix19_En18
  input [18:0] Wgt_8_399, // sfix19_En18
  input [18:0] Wgt_8_400, // sfix19_En18
  input [18:0] Wgt_8_401, // sfix19_En18
  input [18:0] Wgt_8_402, // sfix19_En18
  input [18:0] Wgt_8_403, // sfix19_En18
  input [18:0] Wgt_8_404, // sfix19_En18
  input [18:0] Wgt_8_405, // sfix19_En18
  input [18:0] Wgt_8_406, // sfix19_En18
  input [18:0] Wgt_8_407, // sfix19_En18
  input [18:0] Wgt_8_408, // sfix19_En18
  input [18:0] Wgt_8_409, // sfix19_En18
  input [18:0] Wgt_8_410, // sfix19_En18
  input [18:0] Wgt_8_411, // sfix19_En18
  input [18:0] Wgt_8_412, // sfix19_En18
  input [18:0] Wgt_8_413, // sfix19_En18
  input [18:0] Wgt_8_414, // sfix19_En18
  input [18:0] Wgt_8_415, // sfix19_En18
  input [18:0] Wgt_8_416, // sfix19_En18
  input [18:0] Wgt_8_417, // sfix19_En18
  input [18:0] Wgt_8_418, // sfix19_En18
  input [18:0] Wgt_8_419, // sfix19_En18
  input [18:0] Wgt_8_420, // sfix19_En18
  input [18:0] Wgt_8_421, // sfix19_En18
  input [18:0] Wgt_8_422, // sfix19_En18
  input [18:0] Wgt_8_423, // sfix19_En18
  input [18:0] Wgt_8_424, // sfix19_En18
  input [18:0] Wgt_8_425, // sfix19_En18
  input [18:0] Wgt_8_426, // sfix19_En18
  input [18:0] Wgt_8_427, // sfix19_En18
  input [18:0] Wgt_8_428, // sfix19_En18
  input [18:0] Wgt_8_429, // sfix19_En18
  input [18:0] Wgt_8_430, // sfix19_En18
  input [18:0] Wgt_8_431, // sfix19_En18
  input [18:0] Wgt_8_432, // sfix19_En18
  input [18:0] Wgt_8_433, // sfix19_En18
  input [18:0] Wgt_8_434, // sfix19_En18
  input [18:0] Wgt_8_435, // sfix19_En18
  input [18:0] Wgt_8_436, // sfix19_En18
  input [18:0] Wgt_8_437, // sfix19_En18
  input [18:0] Wgt_8_438, // sfix19_En18
  input [18:0] Wgt_8_439, // sfix19_En18
  input [18:0] Wgt_8_440, // sfix19_En18
  input [18:0] Wgt_8_441, // sfix19_En18
  input [18:0] Wgt_8_442, // sfix19_En18
  input [18:0] Wgt_8_443, // sfix19_En18
  input [18:0] Wgt_8_444, // sfix19_En18
  input [18:0] Wgt_8_445, // sfix19_En18
  input [18:0] Wgt_8_446, // sfix19_En18
  input [18:0] Wgt_8_447, // sfix19_En18
  input [18:0] Wgt_8_448, // sfix19_En18
  input [18:0] Wgt_8_449, // sfix19_En18
  input [18:0] Wgt_8_450, // sfix19_En18
  input [18:0] Wgt_8_451, // sfix19_En18
  input [18:0] Wgt_8_452, // sfix19_En18
  input [18:0] Wgt_8_453, // sfix19_En18
  input [18:0] Wgt_8_454, // sfix19_En18
  input [18:0] Wgt_8_455, // sfix19_En18
  input [18:0] Wgt_8_456, // sfix19_En18
  input [18:0] Wgt_8_457, // sfix19_En18
  input [18:0] Wgt_8_458, // sfix19_En18
  input [18:0] Wgt_8_459, // sfix19_En18
  input [18:0] Wgt_8_460, // sfix19_En18
  input [18:0] Wgt_8_461, // sfix19_En18
  input [18:0] Wgt_8_462, // sfix19_En18
  input [18:0] Wgt_8_463, // sfix19_En18
  input [18:0] Wgt_8_464, // sfix19_En18
  input [18:0] Wgt_8_465, // sfix19_En18
  input [18:0] Wgt_8_466, // sfix19_En18
  input [18:0] Wgt_8_467, // sfix19_En18
  input [18:0] Wgt_8_468, // sfix19_En18
  input [18:0] Wgt_8_469, // sfix19_En18
  input [18:0] Wgt_8_470, // sfix19_En18
  input [18:0] Wgt_8_471, // sfix19_En18
  input [18:0] Wgt_8_472, // sfix19_En18
  input [18:0] Wgt_8_473, // sfix19_En18
  input [18:0] Wgt_8_474, // sfix19_En18
  input [18:0] Wgt_8_475, // sfix19_En18
  input [18:0] Wgt_8_476, // sfix19_En18
  input [18:0] Wgt_8_477, // sfix19_En18
  input [18:0] Wgt_8_478, // sfix19_En18
  input [18:0] Wgt_8_479, // sfix19_En18
  input [18:0] Wgt_8_480, // sfix19_En18
  input [18:0] Wgt_8_481, // sfix19_En18
  input [18:0] Wgt_8_482, // sfix19_En18
  input [18:0] Wgt_8_483, // sfix19_En18
  input [18:0] Wgt_8_484, // sfix19_En18
  input [18:0] Wgt_8_485, // sfix19_En18
  input [18:0] Wgt_8_486, // sfix19_En18
  input [18:0] Wgt_8_487, // sfix19_En18
  input [18:0] Wgt_8_488, // sfix19_En18
  input [18:0] Wgt_8_489, // sfix19_En18
  input [18:0] Wgt_8_490, // sfix19_En18
  input [18:0] Wgt_8_491, // sfix19_En18
  input [18:0] Wgt_8_492, // sfix19_En18
  input [18:0] Wgt_8_493, // sfix19_En18
  input [18:0] Wgt_8_494, // sfix19_En18
  input [18:0] Wgt_8_495, // sfix19_En18
  input [18:0] Wgt_8_496, // sfix19_En18
  input [18:0] Wgt_8_497, // sfix19_En18
  input [18:0] Wgt_8_498, // sfix19_En18
  input [18:0] Wgt_8_499, // sfix19_En18
  input [18:0] Wgt_8_500, // sfix19_En18
  input [18:0] Wgt_8_501, // sfix19_En18
  input [18:0] Wgt_8_502, // sfix19_En18
  input [18:0] Wgt_8_503, // sfix19_En18
  input [18:0] Wgt_8_504, // sfix19_En18
  input [18:0] Wgt_8_505, // sfix19_En18
  input [18:0] Wgt_8_506, // sfix19_En18
  input [18:0] Wgt_8_507, // sfix19_En18
  input [18:0] Wgt_8_508, // sfix19_En18
  input [18:0] Wgt_8_509, // sfix19_En18
  input [18:0] Wgt_8_510, // sfix19_En18
  input [18:0] Wgt_8_511, // sfix19_En18
  input [18:0] Wgt_8_512, // sfix19_En18
  input [18:0] Wgt_8_513, // sfix19_En18
  input [18:0] Wgt_8_514, // sfix19_En18
  input [18:0] Wgt_8_515, // sfix19_En18
  input [18:0] Wgt_8_516, // sfix19_En18
  input [18:0] Wgt_8_517, // sfix19_En18
  input [18:0] Wgt_8_518, // sfix19_En18
  input [18:0] Wgt_8_519, // sfix19_En18
  input [18:0] Wgt_8_520, // sfix19_En18
  input [18:0] Wgt_8_521, // sfix19_En18
  input [18:0] Wgt_8_522, // sfix19_En18
  input [18:0] Wgt_8_523, // sfix19_En18
  input [18:0] Wgt_8_524, // sfix19_En18
  input [18:0] Wgt_8_525, // sfix19_En18
  input [18:0] Wgt_8_526, // sfix19_En18
  input [18:0] Wgt_8_527, // sfix19_En18
  input [18:0] Wgt_8_528, // sfix19_En18
  input [18:0] Wgt_8_529, // sfix19_En18
  input [18:0] Wgt_8_530, // sfix19_En18
  input [18:0] Wgt_8_531, // sfix19_En18
  input [18:0] Wgt_8_532, // sfix19_En18
  input [18:0] Wgt_8_533, // sfix19_En18
  input [18:0] Wgt_8_534, // sfix19_En18
  input [18:0] Wgt_8_535, // sfix19_En18
  input [18:0] Wgt_8_536, // sfix19_En18
  input [18:0] Wgt_8_537, // sfix19_En18
  input [18:0] Wgt_8_538, // sfix19_En18
  input [18:0] Wgt_8_539, // sfix19_En18
  input [18:0] Wgt_8_540, // sfix19_En18
  input [18:0] Wgt_8_541, // sfix19_En18
  input [18:0] Wgt_8_542, // sfix19_En18
  input [18:0] Wgt_8_543, // sfix19_En18
  input [18:0] Wgt_8_544, // sfix19_En18
  input [18:0] Wgt_8_545, // sfix19_En18
  input [18:0] Wgt_8_546, // sfix19_En18
  input [18:0] Wgt_8_547, // sfix19_En18
  input [18:0] Wgt_8_548, // sfix19_En18
  input [18:0] Wgt_8_549, // sfix19_En18
  input [18:0] Wgt_8_550, // sfix19_En18
  input [18:0] Wgt_8_551, // sfix19_En18
  input [18:0] Wgt_8_552, // sfix19_En18
  input [18:0] Wgt_8_553, // sfix19_En18
  input [18:0] Wgt_8_554, // sfix19_En18
  input [18:0] Wgt_8_555, // sfix19_En18
  input [18:0] Wgt_8_556, // sfix19_En18
  input [18:0] Wgt_8_557, // sfix19_En18
  input [18:0] Wgt_8_558, // sfix19_En18
  input [18:0] Wgt_8_559, // sfix19_En18
  input [18:0] Wgt_8_560, // sfix19_En18
  input [18:0] Wgt_8_561, // sfix19_En18
  input [18:0] Wgt_8_562, // sfix19_En18
  input [18:0] Wgt_8_563, // sfix19_En18
  input [18:0] Wgt_8_564, // sfix19_En18
  input [18:0] Wgt_8_565, // sfix19_En18
  input [18:0] Wgt_8_566, // sfix19_En18
  input [18:0] Wgt_8_567, // sfix19_En18
  input [18:0] Wgt_8_568, // sfix19_En18
  input [18:0] Wgt_8_569, // sfix19_En18
  input [18:0] Wgt_8_570, // sfix19_En18
  input [18:0] Wgt_8_571, // sfix19_En18
  input [18:0] Wgt_8_572, // sfix19_En18
  input [18:0] Wgt_8_573, // sfix19_En18
  input [18:0] Wgt_8_574, // sfix19_En18
  input [18:0] Wgt_8_575, // sfix19_En18
  input [18:0] Wgt_8_576, // sfix19_En18
  input [18:0] Wgt_8_577, // sfix19_En18
  input [18:0] Wgt_8_578, // sfix19_En18
  input [18:0] Wgt_8_579, // sfix19_En18
  input [18:0] Wgt_8_580, // sfix19_En18
  input [18:0] Wgt_8_581, // sfix19_En18
  input [18:0] Wgt_8_582, // sfix19_En18
  input [18:0] Wgt_8_583, // sfix19_En18
  input [18:0] Wgt_8_584, // sfix19_En18
  input [18:0] Wgt_8_585, // sfix19_En18
  input [18:0] Wgt_8_586, // sfix19_En18
  input [18:0] Wgt_8_587, // sfix19_En18
  input [18:0] Wgt_8_588, // sfix19_En18
  input [18:0] Wgt_8_589, // sfix19_En18
  input [18:0] Wgt_8_590, // sfix19_En18
  input [18:0] Wgt_8_591, // sfix19_En18
  input [18:0] Wgt_8_592, // sfix19_En18
  input [18:0] Wgt_8_593, // sfix19_En18
  input [18:0] Wgt_8_594, // sfix19_En18
  input [18:0] Wgt_8_595, // sfix19_En18
  input [18:0] Wgt_8_596, // sfix19_En18
  input [18:0] Wgt_8_597, // sfix19_En18
  input [18:0] Wgt_8_598, // sfix19_En18
  input [18:0] Wgt_8_599, // sfix19_En18
  input [18:0] Wgt_8_600, // sfix19_En18
  input [18:0] Wgt_8_601, // sfix19_En18
  input [18:0] Wgt_8_602, // sfix19_En18
  input [18:0] Wgt_8_603, // sfix19_En18
  input [18:0] Wgt_8_604, // sfix19_En18
  input [18:0] Wgt_8_605, // sfix19_En18
  input [18:0] Wgt_8_606, // sfix19_En18
  input [18:0] Wgt_8_607, // sfix19_En18
  input [18:0] Wgt_8_608, // sfix19_En18
  input [18:0] Wgt_8_609, // sfix19_En18
  input [18:0] Wgt_8_610, // sfix19_En18
  input [18:0] Wgt_8_611, // sfix19_En18
  input [18:0] Wgt_8_612, // sfix19_En18
  input [18:0] Wgt_8_613, // sfix19_En18
  input [18:0] Wgt_8_614, // sfix19_En18
  input [18:0] Wgt_8_615, // sfix19_En18
  input [18:0] Wgt_8_616, // sfix19_En18
  input [18:0] Wgt_8_617, // sfix19_En18
  input [18:0] Wgt_8_618, // sfix19_En18
  input [18:0] Wgt_8_619, // sfix19_En18
  input [18:0] Wgt_8_620, // sfix19_En18
  input [18:0] Wgt_8_621, // sfix19_En18
  input [18:0] Wgt_8_622, // sfix19_En18
  input [18:0] Wgt_8_623, // sfix19_En18
  input [18:0] Wgt_8_624, // sfix19_En18
  input [18:0] Wgt_8_625, // sfix19_En18
  input [18:0] Wgt_8_626, // sfix19_En18
  input [18:0] Wgt_8_627, // sfix19_En18
  input [18:0] Wgt_8_628, // sfix19_En18
  input [18:0] Wgt_8_629, // sfix19_En18
  input [18:0] Wgt_8_630, // sfix19_En18
  input [18:0] Wgt_8_631, // sfix19_En18
  input [18:0] Wgt_8_632, // sfix19_En18
  input [18:0] Wgt_8_633, // sfix19_En18
  input [18:0] Wgt_8_634, // sfix19_En18
  input [18:0] Wgt_8_635, // sfix19_En18
  input [18:0] Wgt_8_636, // sfix19_En18
  input [18:0] Wgt_8_637, // sfix19_En18
  input [18:0] Wgt_8_638, // sfix19_En18
  input [18:0] Wgt_8_639, // sfix19_En18
  input [18:0] Wgt_8_640, // sfix19_En18
  input [18:0] Wgt_8_641, // sfix19_En18
  input [18:0] Wgt_8_642, // sfix19_En18
  input [18:0] Wgt_8_643, // sfix19_En18
  input [18:0] Wgt_8_644, // sfix19_En18
  input [18:0] Wgt_8_645, // sfix19_En18
  input [18:0] Wgt_8_646, // sfix19_En18
  input [18:0] Wgt_8_647, // sfix19_En18
  input [18:0] Wgt_8_648, // sfix19_En18
  input [18:0] Wgt_8_649, // sfix19_En18
  input [18:0] Wgt_8_650, // sfix19_En18
  input [18:0] Wgt_8_651, // sfix19_En18
  input [18:0] Wgt_8_652, // sfix19_En18
  input [18:0] Wgt_8_653, // sfix19_En18
  input [18:0] Wgt_8_654, // sfix19_En18
  input [18:0] Wgt_8_655, // sfix19_En18
  input [18:0] Wgt_8_656, // sfix19_En18
  input [18:0] Wgt_8_657, // sfix19_En18
  input [18:0] Wgt_8_658, // sfix19_En18
  input [18:0] Wgt_8_659, // sfix19_En18
  input [18:0] Wgt_8_660, // sfix19_En18
  input [18:0] Wgt_8_661, // sfix19_En18
  input [18:0] Wgt_8_662, // sfix19_En18
  input [18:0] Wgt_8_663, // sfix19_En18
  input [18:0] Wgt_8_664, // sfix19_En18
  input [18:0] Wgt_8_665, // sfix19_En18
  input [18:0] Wgt_8_666, // sfix19_En18
  input [18:0] Wgt_8_667, // sfix19_En18
  input [18:0] Wgt_8_668, // sfix19_En18
  input [18:0] Wgt_8_669, // sfix19_En18
  input [18:0] Wgt_8_670, // sfix19_En18
  input [18:0] Wgt_8_671, // sfix19_En18
  input [18:0] Wgt_8_672, // sfix19_En18
  input [18:0] Wgt_8_673, // sfix19_En18
  input [18:0] Wgt_8_674, // sfix19_En18
  input [18:0] Wgt_8_675, // sfix19_En18
  input [18:0] Wgt_8_676, // sfix19_En18
  input [18:0] Wgt_8_677, // sfix19_En18
  input [18:0] Wgt_8_678, // sfix19_En18
  input [18:0] Wgt_8_679, // sfix19_En18
  input [18:0] Wgt_8_680, // sfix19_En18
  input [18:0] Wgt_8_681, // sfix19_En18
  input [18:0] Wgt_8_682, // sfix19_En18
  input [18:0] Wgt_8_683, // sfix19_En18
  input [18:0] Wgt_8_684, // sfix19_En18
  input [18:0] Wgt_8_685, // sfix19_En18
  input [18:0] Wgt_8_686, // sfix19_En18
  input [18:0] Wgt_8_687, // sfix19_En18
  input [18:0] Wgt_8_688, // sfix19_En18
  input [18:0] Wgt_8_689, // sfix19_En18
  input [18:0] Wgt_8_690, // sfix19_En18
  input [18:0] Wgt_8_691, // sfix19_En18
  input [18:0] Wgt_8_692, // sfix19_En18
  input [18:0] Wgt_8_693, // sfix19_En18
  input [18:0] Wgt_8_694, // sfix19_En18
  input [18:0] Wgt_8_695, // sfix19_En18
  input [18:0] Wgt_8_696, // sfix19_En18
  input [18:0] Wgt_8_697, // sfix19_En18
  input [18:0] Wgt_8_698, // sfix19_En18
  input [18:0] Wgt_8_699, // sfix19_En18
  input [18:0] Wgt_8_700, // sfix19_En18
  input [18:0] Wgt_8_701, // sfix19_En18
  input [18:0] Wgt_8_702, // sfix19_En18
  input [18:0] Wgt_8_703, // sfix19_En18
  input [18:0] Wgt_8_704, // sfix19_En18
  input [18:0] Wgt_8_705, // sfix19_En18
  input [18:0] Wgt_8_706, // sfix19_En18
  input [18:0] Wgt_8_707, // sfix19_En18
  input [18:0] Wgt_8_708, // sfix19_En18
  input [18:0] Wgt_8_709, // sfix19_En18
  input [18:0] Wgt_8_710, // sfix19_En18
  input [18:0] Wgt_8_711, // sfix19_En18
  input [18:0] Wgt_8_712, // sfix19_En18
  input [18:0] Wgt_8_713, // sfix19_En18
  input [18:0] Wgt_8_714, // sfix19_En18
  input [18:0] Wgt_8_715, // sfix19_En18
  input [18:0] Wgt_8_716, // sfix19_En18
  input [18:0] Wgt_8_717, // sfix19_En18
  input [18:0] Wgt_8_718, // sfix19_En18
  input [18:0] Wgt_8_719, // sfix19_En18
  input [18:0] Wgt_8_720, // sfix19_En18
  input [18:0] Wgt_8_721, // sfix19_En18
  input [18:0] Wgt_8_722, // sfix19_En18
  input [18:0] Wgt_8_723, // sfix19_En18
  input [18:0] Wgt_8_724, // sfix19_En18
  input [18:0] Wgt_8_725, // sfix19_En18
  input [18:0] Wgt_8_726, // sfix19_En18
  input [18:0] Wgt_8_727, // sfix19_En18
  input [18:0] Wgt_8_728, // sfix19_En18
  input [18:0] Wgt_8_729, // sfix19_En18
  input [18:0] Wgt_8_730, // sfix19_En18
  input [18:0] Wgt_8_731, // sfix19_En18
  input [18:0] Wgt_8_732, // sfix19_En18
  input [18:0] Wgt_8_733, // sfix19_En18
  input [18:0] Wgt_8_734, // sfix19_En18
  input [18:0] Wgt_8_735, // sfix19_En18
  input [18:0] Wgt_8_736, // sfix19_En18
  input [18:0] Wgt_8_737, // sfix19_En18
  input [18:0] Wgt_8_738, // sfix19_En18
  input [18:0] Wgt_8_739, // sfix19_En18
  input [18:0] Wgt_8_740, // sfix19_En18
  input [18:0] Wgt_8_741, // sfix19_En18
  input [18:0] Wgt_8_742, // sfix19_En18
  input [18:0] Wgt_8_743, // sfix19_En18
  input [18:0] Wgt_8_744, // sfix19_En18
  input [18:0] Wgt_8_745, // sfix19_En18
  input [18:0] Wgt_8_746, // sfix19_En18
  input [18:0] Wgt_8_747, // sfix19_En18
  input [18:0] Wgt_8_748, // sfix19_En18
  input [18:0] Wgt_8_749, // sfix19_En18
  input [18:0] Wgt_8_750, // sfix19_En18
  input [18:0] Wgt_8_751, // sfix19_En18
  input [18:0] Wgt_8_752, // sfix19_En18
  input [18:0] Wgt_8_753, // sfix19_En18
  input [18:0] Wgt_8_754, // sfix19_En18
  input [18:0] Wgt_8_755, // sfix19_En18
  input [18:0] Wgt_8_756, // sfix19_En18
  input [18:0] Wgt_8_757, // sfix19_En18
  input [18:0] Wgt_8_758, // sfix19_En18
  input [18:0] Wgt_8_759, // sfix19_En18
  input [18:0] Wgt_8_760, // sfix19_En18
  input [18:0] Wgt_8_761, // sfix19_En18
  input [18:0] Wgt_8_762, // sfix19_En18
  input [18:0] Wgt_8_763, // sfix19_En18
  input [18:0] Wgt_8_764, // sfix19_En18
  input [18:0] Wgt_8_765, // sfix19_En18
  input [18:0] Wgt_8_766, // sfix19_En18
  input [18:0] Wgt_8_767, // sfix19_En18
  input [18:0] Wgt_8_768, // sfix19_En18
  input [18:0] Wgt_8_769, // sfix19_En18
  input [18:0] Wgt_8_770, // sfix19_En18
  input [18:0] Wgt_8_771, // sfix19_En18
  input [18:0] Wgt_8_772, // sfix19_En18
  input [18:0] Wgt_8_773, // sfix19_En18
  input [18:0] Wgt_8_774, // sfix19_En18
  input [18:0] Wgt_8_775, // sfix19_En18
  input [18:0] Wgt_8_776, // sfix19_En18
  input [18:0] Wgt_8_777, // sfix19_En18
  input [18:0] Wgt_8_778, // sfix19_En18
  input [18:0] Wgt_8_779, // sfix19_En18
  input [18:0] Wgt_8_780, // sfix19_En18
  input [18:0] Wgt_8_781, // sfix19_En18
  input [18:0] Wgt_8_782, // sfix19_En18
  input [18:0] Wgt_8_783, // sfix19_En18
  input [18:0] Wgt_8_784, // sfix19_En18
  input [18:0] Wgt_9_0, // sfix19_En18
  input [18:0] Wgt_9_1, // sfix19_En18
  input [18:0] Wgt_9_2, // sfix19_En18
  input [18:0] Wgt_9_3, // sfix19_En18
  input [18:0] Wgt_9_4, // sfix19_En18
  input [18:0] Wgt_9_5, // sfix19_En18
  input [18:0] Wgt_9_6, // sfix19_En18
  input [18:0] Wgt_9_7, // sfix19_En18
  input [18:0] Wgt_9_8, // sfix19_En18
  input [18:0] Wgt_9_9, // sfix19_En18
  input [18:0] Wgt_9_10, // sfix19_En18
  input [18:0] Wgt_9_11, // sfix19_En18
  input [18:0] Wgt_9_12, // sfix19_En18
  input [18:0] Wgt_9_13, // sfix19_En18
  input [18:0] Wgt_9_14, // sfix19_En18
  input [18:0] Wgt_9_15, // sfix19_En18
  input [18:0] Wgt_9_16, // sfix19_En18
  input [18:0] Wgt_9_17, // sfix19_En18
  input [18:0] Wgt_9_18, // sfix19_En18
  input [18:0] Wgt_9_19, // sfix19_En18
  input [18:0] Wgt_9_20, // sfix19_En18
  input [18:0] Wgt_9_21, // sfix19_En18
  input [18:0] Wgt_9_22, // sfix19_En18
  input [18:0] Wgt_9_23, // sfix19_En18
  input [18:0] Wgt_9_24, // sfix19_En18
  input [18:0] Wgt_9_25, // sfix19_En18
  input [18:0] Wgt_9_26, // sfix19_En18
  input [18:0] Wgt_9_27, // sfix19_En18
  input [18:0] Wgt_9_28, // sfix19_En18
  input [18:0] Wgt_9_29, // sfix19_En18
  input [18:0] Wgt_9_30, // sfix19_En18
  input [18:0] Wgt_9_31, // sfix19_En18
  input [18:0] Wgt_9_32, // sfix19_En18
  input [18:0] Wgt_9_33, // sfix19_En18
  input [18:0] Wgt_9_34, // sfix19_En18
  input [18:0] Wgt_9_35, // sfix19_En18
  input [18:0] Wgt_9_36, // sfix19_En18
  input [18:0] Wgt_9_37, // sfix19_En18
  input [18:0] Wgt_9_38, // sfix19_En18
  input [18:0] Wgt_9_39, // sfix19_En18
  input [18:0] Wgt_9_40, // sfix19_En18
  input [18:0] Wgt_9_41, // sfix19_En18
  input [18:0] Wgt_9_42, // sfix19_En18
  input [18:0] Wgt_9_43, // sfix19_En18
  input [18:0] Wgt_9_44, // sfix19_En18
  input [18:0] Wgt_9_45, // sfix19_En18
  input [18:0] Wgt_9_46, // sfix19_En18
  input [18:0] Wgt_9_47, // sfix19_En18
  input [18:0] Wgt_9_48, // sfix19_En18
  input [18:0] Wgt_9_49, // sfix19_En18
  input [18:0] Wgt_9_50, // sfix19_En18
  input [18:0] Wgt_9_51, // sfix19_En18
  input [18:0] Wgt_9_52, // sfix19_En18
  input [18:0] Wgt_9_53, // sfix19_En18
  input [18:0] Wgt_9_54, // sfix19_En18
  input [18:0] Wgt_9_55, // sfix19_En18
  input [18:0] Wgt_9_56, // sfix19_En18
  input [18:0] Wgt_9_57, // sfix19_En18
  input [18:0] Wgt_9_58, // sfix19_En18
  input [18:0] Wgt_9_59, // sfix19_En18
  input [18:0] Wgt_9_60, // sfix19_En18
  input [18:0] Wgt_9_61, // sfix19_En18
  input [18:0] Wgt_9_62, // sfix19_En18
  input [18:0] Wgt_9_63, // sfix19_En18
  input [18:0] Wgt_9_64, // sfix19_En18
  input [18:0] Wgt_9_65, // sfix19_En18
  input [18:0] Wgt_9_66, // sfix19_En18
  input [18:0] Wgt_9_67, // sfix19_En18
  input [18:0] Wgt_9_68, // sfix19_En18
  input [18:0] Wgt_9_69, // sfix19_En18
  input [18:0] Wgt_9_70, // sfix19_En18
  input [18:0] Wgt_9_71, // sfix19_En18
  input [18:0] Wgt_9_72, // sfix19_En18
  input [18:0] Wgt_9_73, // sfix19_En18
  input [18:0] Wgt_9_74, // sfix19_En18
  input [18:0] Wgt_9_75, // sfix19_En18
  input [18:0] Wgt_9_76, // sfix19_En18
  input [18:0] Wgt_9_77, // sfix19_En18
  input [18:0] Wgt_9_78, // sfix19_En18
  input [18:0] Wgt_9_79, // sfix19_En18
  input [18:0] Wgt_9_80, // sfix19_En18
  input [18:0] Wgt_9_81, // sfix19_En18
  input [18:0] Wgt_9_82, // sfix19_En18
  input [18:0] Wgt_9_83, // sfix19_En18
  input [18:0] Wgt_9_84, // sfix19_En18
  input [18:0] Wgt_9_85, // sfix19_En18
  input [18:0] Wgt_9_86, // sfix19_En18
  input [18:0] Wgt_9_87, // sfix19_En18
  input [18:0] Wgt_9_88, // sfix19_En18
  input [18:0] Wgt_9_89, // sfix19_En18
  input [18:0] Wgt_9_90, // sfix19_En18
  input [18:0] Wgt_9_91, // sfix19_En18
  input [18:0] Wgt_9_92, // sfix19_En18
  input [18:0] Wgt_9_93, // sfix19_En18
  input [18:0] Wgt_9_94, // sfix19_En18
  input [18:0] Wgt_9_95, // sfix19_En18
  input [18:0] Wgt_9_96, // sfix19_En18
  input [18:0] Wgt_9_97, // sfix19_En18
  input [18:0] Wgt_9_98, // sfix19_En18
  input [18:0] Wgt_9_99, // sfix19_En18
  input [18:0] Wgt_9_100, // sfix19_En18
  input [18:0] Wgt_9_101, // sfix19_En18
  input [18:0] Wgt_9_102, // sfix19_En18
  input [18:0] Wgt_9_103, // sfix19_En18
  input [18:0] Wgt_9_104, // sfix19_En18
  input [18:0] Wgt_9_105, // sfix19_En18
  input [18:0] Wgt_9_106, // sfix19_En18
  input [18:0] Wgt_9_107, // sfix19_En18
  input [18:0] Wgt_9_108, // sfix19_En18
  input [18:0] Wgt_9_109, // sfix19_En18
  input [18:0] Wgt_9_110, // sfix19_En18
  input [18:0] Wgt_9_111, // sfix19_En18
  input [18:0] Wgt_9_112, // sfix19_En18
  input [18:0] Wgt_9_113, // sfix19_En18
  input [18:0] Wgt_9_114, // sfix19_En18
  input [18:0] Wgt_9_115, // sfix19_En18
  input [18:0] Wgt_9_116, // sfix19_En18
  input [18:0] Wgt_9_117, // sfix19_En18
  input [18:0] Wgt_9_118, // sfix19_En18
  input [18:0] Wgt_9_119, // sfix19_En18
  input [18:0] Wgt_9_120, // sfix19_En18
  input [18:0] Wgt_9_121, // sfix19_En18
  input [18:0] Wgt_9_122, // sfix19_En18
  input [18:0] Wgt_9_123, // sfix19_En18
  input [18:0] Wgt_9_124, // sfix19_En18
  input [18:0] Wgt_9_125, // sfix19_En18
  input [18:0] Wgt_9_126, // sfix19_En18
  input [18:0] Wgt_9_127, // sfix19_En18
  input [18:0] Wgt_9_128, // sfix19_En18
  input [18:0] Wgt_9_129, // sfix19_En18
  input [18:0] Wgt_9_130, // sfix19_En18
  input [18:0] Wgt_9_131, // sfix19_En18
  input [18:0] Wgt_9_132, // sfix19_En18
  input [18:0] Wgt_9_133, // sfix19_En18
  input [18:0] Wgt_9_134, // sfix19_En18
  input [18:0] Wgt_9_135, // sfix19_En18
  input [18:0] Wgt_9_136, // sfix19_En18
  input [18:0] Wgt_9_137, // sfix19_En18
  input [18:0] Wgt_9_138, // sfix19_En18
  input [18:0] Wgt_9_139, // sfix19_En18
  input [18:0] Wgt_9_140, // sfix19_En18
  input [18:0] Wgt_9_141, // sfix19_En18
  input [18:0] Wgt_9_142, // sfix19_En18
  input [18:0] Wgt_9_143, // sfix19_En18
  input [18:0] Wgt_9_144, // sfix19_En18
  input [18:0] Wgt_9_145, // sfix19_En18
  input [18:0] Wgt_9_146, // sfix19_En18
  input [18:0] Wgt_9_147, // sfix19_En18
  input [18:0] Wgt_9_148, // sfix19_En18
  input [18:0] Wgt_9_149, // sfix19_En18
  input [18:0] Wgt_9_150, // sfix19_En18
  input [18:0] Wgt_9_151, // sfix19_En18
  input [18:0] Wgt_9_152, // sfix19_En18
  input [18:0] Wgt_9_153, // sfix19_En18
  input [18:0] Wgt_9_154, // sfix19_En18
  input [18:0] Wgt_9_155, // sfix19_En18
  input [18:0] Wgt_9_156, // sfix19_En18
  input [18:0] Wgt_9_157, // sfix19_En18
  input [18:0] Wgt_9_158, // sfix19_En18
  input [18:0] Wgt_9_159, // sfix19_En18
  input [18:0] Wgt_9_160, // sfix19_En18
  input [18:0] Wgt_9_161, // sfix19_En18
  input [18:0] Wgt_9_162, // sfix19_En18
  input [18:0] Wgt_9_163, // sfix19_En18
  input [18:0] Wgt_9_164, // sfix19_En18
  input [18:0] Wgt_9_165, // sfix19_En18
  input [18:0] Wgt_9_166, // sfix19_En18
  input [18:0] Wgt_9_167, // sfix19_En18
  input [18:0] Wgt_9_168, // sfix19_En18
  input [18:0] Wgt_9_169, // sfix19_En18
  input [18:0] Wgt_9_170, // sfix19_En18
  input [18:0] Wgt_9_171, // sfix19_En18
  input [18:0] Wgt_9_172, // sfix19_En18
  input [18:0] Wgt_9_173, // sfix19_En18
  input [18:0] Wgt_9_174, // sfix19_En18
  input [18:0] Wgt_9_175, // sfix19_En18
  input [18:0] Wgt_9_176, // sfix19_En18
  input [18:0] Wgt_9_177, // sfix19_En18
  input [18:0] Wgt_9_178, // sfix19_En18
  input [18:0] Wgt_9_179, // sfix19_En18
  input [18:0] Wgt_9_180, // sfix19_En18
  input [18:0] Wgt_9_181, // sfix19_En18
  input [18:0] Wgt_9_182, // sfix19_En18
  input [18:0] Wgt_9_183, // sfix19_En18
  input [18:0] Wgt_9_184, // sfix19_En18
  input [18:0] Wgt_9_185, // sfix19_En18
  input [18:0] Wgt_9_186, // sfix19_En18
  input [18:0] Wgt_9_187, // sfix19_En18
  input [18:0] Wgt_9_188, // sfix19_En18
  input [18:0] Wgt_9_189, // sfix19_En18
  input [18:0] Wgt_9_190, // sfix19_En18
  input [18:0] Wgt_9_191, // sfix19_En18
  input [18:0] Wgt_9_192, // sfix19_En18
  input [18:0] Wgt_9_193, // sfix19_En18
  input [18:0] Wgt_9_194, // sfix19_En18
  input [18:0] Wgt_9_195, // sfix19_En18
  input [18:0] Wgt_9_196, // sfix19_En18
  input [18:0] Wgt_9_197, // sfix19_En18
  input [18:0] Wgt_9_198, // sfix19_En18
  input [18:0] Wgt_9_199, // sfix19_En18
  input [18:0] Wgt_9_200, // sfix19_En18
  input [18:0] Wgt_9_201, // sfix19_En18
  input [18:0] Wgt_9_202, // sfix19_En18
  input [18:0] Wgt_9_203, // sfix19_En18
  input [18:0] Wgt_9_204, // sfix19_En18
  input [18:0] Wgt_9_205, // sfix19_En18
  input [18:0] Wgt_9_206, // sfix19_En18
  input [18:0] Wgt_9_207, // sfix19_En18
  input [18:0] Wgt_9_208, // sfix19_En18
  input [18:0] Wgt_9_209, // sfix19_En18
  input [18:0] Wgt_9_210, // sfix19_En18
  input [18:0] Wgt_9_211, // sfix19_En18
  input [18:0] Wgt_9_212, // sfix19_En18
  input [18:0] Wgt_9_213, // sfix19_En18
  input [18:0] Wgt_9_214, // sfix19_En18
  input [18:0] Wgt_9_215, // sfix19_En18
  input [18:0] Wgt_9_216, // sfix19_En18
  input [18:0] Wgt_9_217, // sfix19_En18
  input [18:0] Wgt_9_218, // sfix19_En18
  input [18:0] Wgt_9_219, // sfix19_En18
  input [18:0] Wgt_9_220, // sfix19_En18
  input [18:0] Wgt_9_221, // sfix19_En18
  input [18:0] Wgt_9_222, // sfix19_En18
  input [18:0] Wgt_9_223, // sfix19_En18
  input [18:0] Wgt_9_224, // sfix19_En18
  input [18:0] Wgt_9_225, // sfix19_En18
  input [18:0] Wgt_9_226, // sfix19_En18
  input [18:0] Wgt_9_227, // sfix19_En18
  input [18:0] Wgt_9_228, // sfix19_En18
  input [18:0] Wgt_9_229, // sfix19_En18
  input [18:0] Wgt_9_230, // sfix19_En18
  input [18:0] Wgt_9_231, // sfix19_En18
  input [18:0] Wgt_9_232, // sfix19_En18
  input [18:0] Wgt_9_233, // sfix19_En18
  input [18:0] Wgt_9_234, // sfix19_En18
  input [18:0] Wgt_9_235, // sfix19_En18
  input [18:0] Wgt_9_236, // sfix19_En18
  input [18:0] Wgt_9_237, // sfix19_En18
  input [18:0] Wgt_9_238, // sfix19_En18
  input [18:0] Wgt_9_239, // sfix19_En18
  input [18:0] Wgt_9_240, // sfix19_En18
  input [18:0] Wgt_9_241, // sfix19_En18
  input [18:0] Wgt_9_242, // sfix19_En18
  input [18:0] Wgt_9_243, // sfix19_En18
  input [18:0] Wgt_9_244, // sfix19_En18
  input [18:0] Wgt_9_245, // sfix19_En18
  input [18:0] Wgt_9_246, // sfix19_En18
  input [18:0] Wgt_9_247, // sfix19_En18
  input [18:0] Wgt_9_248, // sfix19_En18
  input [18:0] Wgt_9_249, // sfix19_En18
  input [18:0] Wgt_9_250, // sfix19_En18
  input [18:0] Wgt_9_251, // sfix19_En18
  input [18:0] Wgt_9_252, // sfix19_En18
  input [18:0] Wgt_9_253, // sfix19_En18
  input [18:0] Wgt_9_254, // sfix19_En18
  input [18:0] Wgt_9_255, // sfix19_En18
  input [18:0] Wgt_9_256, // sfix19_En18
  input [18:0] Wgt_9_257, // sfix19_En18
  input [18:0] Wgt_9_258, // sfix19_En18
  input [18:0] Wgt_9_259, // sfix19_En18
  input [18:0] Wgt_9_260, // sfix19_En18
  input [18:0] Wgt_9_261, // sfix19_En18
  input [18:0] Wgt_9_262, // sfix19_En18
  input [18:0] Wgt_9_263, // sfix19_En18
  input [18:0] Wgt_9_264, // sfix19_En18
  input [18:0] Wgt_9_265, // sfix19_En18
  input [18:0] Wgt_9_266, // sfix19_En18
  input [18:0] Wgt_9_267, // sfix19_En18
  input [18:0] Wgt_9_268, // sfix19_En18
  input [18:0] Wgt_9_269, // sfix19_En18
  input [18:0] Wgt_9_270, // sfix19_En18
  input [18:0] Wgt_9_271, // sfix19_En18
  input [18:0] Wgt_9_272, // sfix19_En18
  input [18:0] Wgt_9_273, // sfix19_En18
  input [18:0] Wgt_9_274, // sfix19_En18
  input [18:0] Wgt_9_275, // sfix19_En18
  input [18:0] Wgt_9_276, // sfix19_En18
  input [18:0] Wgt_9_277, // sfix19_En18
  input [18:0] Wgt_9_278, // sfix19_En18
  input [18:0] Wgt_9_279, // sfix19_En18
  input [18:0] Wgt_9_280, // sfix19_En18
  input [18:0] Wgt_9_281, // sfix19_En18
  input [18:0] Wgt_9_282, // sfix19_En18
  input [18:0] Wgt_9_283, // sfix19_En18
  input [18:0] Wgt_9_284, // sfix19_En18
  input [18:0] Wgt_9_285, // sfix19_En18
  input [18:0] Wgt_9_286, // sfix19_En18
  input [18:0] Wgt_9_287, // sfix19_En18
  input [18:0] Wgt_9_288, // sfix19_En18
  input [18:0] Wgt_9_289, // sfix19_En18
  input [18:0] Wgt_9_290, // sfix19_En18
  input [18:0] Wgt_9_291, // sfix19_En18
  input [18:0] Wgt_9_292, // sfix19_En18
  input [18:0] Wgt_9_293, // sfix19_En18
  input [18:0] Wgt_9_294, // sfix19_En18
  input [18:0] Wgt_9_295, // sfix19_En18
  input [18:0] Wgt_9_296, // sfix19_En18
  input [18:0] Wgt_9_297, // sfix19_En18
  input [18:0] Wgt_9_298, // sfix19_En18
  input [18:0] Wgt_9_299, // sfix19_En18
  input [18:0] Wgt_9_300, // sfix19_En18
  input [18:0] Wgt_9_301, // sfix19_En18
  input [18:0] Wgt_9_302, // sfix19_En18
  input [18:0] Wgt_9_303, // sfix19_En18
  input [18:0] Wgt_9_304, // sfix19_En18
  input [18:0] Wgt_9_305, // sfix19_En18
  input [18:0] Wgt_9_306, // sfix19_En18
  input [18:0] Wgt_9_307, // sfix19_En18
  input [18:0] Wgt_9_308, // sfix19_En18
  input [18:0] Wgt_9_309, // sfix19_En18
  input [18:0] Wgt_9_310, // sfix19_En18
  input [18:0] Wgt_9_311, // sfix19_En18
  input [18:0] Wgt_9_312, // sfix19_En18
  input [18:0] Wgt_9_313, // sfix19_En18
  input [18:0] Wgt_9_314, // sfix19_En18
  input [18:0] Wgt_9_315, // sfix19_En18
  input [18:0] Wgt_9_316, // sfix19_En18
  input [18:0] Wgt_9_317, // sfix19_En18
  input [18:0] Wgt_9_318, // sfix19_En18
  input [18:0] Wgt_9_319, // sfix19_En18
  input [18:0] Wgt_9_320, // sfix19_En18
  input [18:0] Wgt_9_321, // sfix19_En18
  input [18:0] Wgt_9_322, // sfix19_En18
  input [18:0] Wgt_9_323, // sfix19_En18
  input [18:0] Wgt_9_324, // sfix19_En18
  input [18:0] Wgt_9_325, // sfix19_En18
  input [18:0] Wgt_9_326, // sfix19_En18
  input [18:0] Wgt_9_327, // sfix19_En18
  input [18:0] Wgt_9_328, // sfix19_En18
  input [18:0] Wgt_9_329, // sfix19_En18
  input [18:0] Wgt_9_330, // sfix19_En18
  input [18:0] Wgt_9_331, // sfix19_En18
  input [18:0] Wgt_9_332, // sfix19_En18
  input [18:0] Wgt_9_333, // sfix19_En18
  input [18:0] Wgt_9_334, // sfix19_En18
  input [18:0] Wgt_9_335, // sfix19_En18
  input [18:0] Wgt_9_336, // sfix19_En18
  input [18:0] Wgt_9_337, // sfix19_En18
  input [18:0] Wgt_9_338, // sfix19_En18
  input [18:0] Wgt_9_339, // sfix19_En18
  input [18:0] Wgt_9_340, // sfix19_En18
  input [18:0] Wgt_9_341, // sfix19_En18
  input [18:0] Wgt_9_342, // sfix19_En18
  input [18:0] Wgt_9_343, // sfix19_En18
  input [18:0] Wgt_9_344, // sfix19_En18
  input [18:0] Wgt_9_345, // sfix19_En18
  input [18:0] Wgt_9_346, // sfix19_En18
  input [18:0] Wgt_9_347, // sfix19_En18
  input [18:0] Wgt_9_348, // sfix19_En18
  input [18:0] Wgt_9_349, // sfix19_En18
  input [18:0] Wgt_9_350, // sfix19_En18
  input [18:0] Wgt_9_351, // sfix19_En18
  input [18:0] Wgt_9_352, // sfix19_En18
  input [18:0] Wgt_9_353, // sfix19_En18
  input [18:0] Wgt_9_354, // sfix19_En18
  input [18:0] Wgt_9_355, // sfix19_En18
  input [18:0] Wgt_9_356, // sfix19_En18
  input [18:0] Wgt_9_357, // sfix19_En18
  input [18:0] Wgt_9_358, // sfix19_En18
  input [18:0] Wgt_9_359, // sfix19_En18
  input [18:0] Wgt_9_360, // sfix19_En18
  input [18:0] Wgt_9_361, // sfix19_En18
  input [18:0] Wgt_9_362, // sfix19_En18
  input [18:0] Wgt_9_363, // sfix19_En18
  input [18:0] Wgt_9_364, // sfix19_En18
  input [18:0] Wgt_9_365, // sfix19_En18
  input [18:0] Wgt_9_366, // sfix19_En18
  input [18:0] Wgt_9_367, // sfix19_En18
  input [18:0] Wgt_9_368, // sfix19_En18
  input [18:0] Wgt_9_369, // sfix19_En18
  input [18:0] Wgt_9_370, // sfix19_En18
  input [18:0] Wgt_9_371, // sfix19_En18
  input [18:0] Wgt_9_372, // sfix19_En18
  input [18:0] Wgt_9_373, // sfix19_En18
  input [18:0] Wgt_9_374, // sfix19_En18
  input [18:0] Wgt_9_375, // sfix19_En18
  input [18:0] Wgt_9_376, // sfix19_En18
  input [18:0] Wgt_9_377, // sfix19_En18
  input [18:0] Wgt_9_378, // sfix19_En18
  input [18:0] Wgt_9_379, // sfix19_En18
  input [18:0] Wgt_9_380, // sfix19_En18
  input [18:0] Wgt_9_381, // sfix19_En18
  input [18:0] Wgt_9_382, // sfix19_En18
  input [18:0] Wgt_9_383, // sfix19_En18
  input [18:0] Wgt_9_384, // sfix19_En18
  input [18:0] Wgt_9_385, // sfix19_En18
  input [18:0] Wgt_9_386, // sfix19_En18
  input [18:0] Wgt_9_387, // sfix19_En18
  input [18:0] Wgt_9_388, // sfix19_En18
  input [18:0] Wgt_9_389, // sfix19_En18
  input [18:0] Wgt_9_390, // sfix19_En18
  input [18:0] Wgt_9_391, // sfix19_En18
  input [18:0] Wgt_9_392, // sfix19_En18
  input [18:0] Wgt_9_393, // sfix19_En18
  input [18:0] Wgt_9_394, // sfix19_En18
  input [18:0] Wgt_9_395, // sfix19_En18
  input [18:0] Wgt_9_396, // sfix19_En18
  input [18:0] Wgt_9_397, // sfix19_En18
  input [18:0] Wgt_9_398, // sfix19_En18
  input [18:0] Wgt_9_399, // sfix19_En18
  input [18:0] Wgt_9_400, // sfix19_En18
  input [18:0] Wgt_9_401, // sfix19_En18
  input [18:0] Wgt_9_402, // sfix19_En18
  input [18:0] Wgt_9_403, // sfix19_En18
  input [18:0] Wgt_9_404, // sfix19_En18
  input [18:0] Wgt_9_405, // sfix19_En18
  input [18:0] Wgt_9_406, // sfix19_En18
  input [18:0] Wgt_9_407, // sfix19_En18
  input [18:0] Wgt_9_408, // sfix19_En18
  input [18:0] Wgt_9_409, // sfix19_En18
  input [18:0] Wgt_9_410, // sfix19_En18
  input [18:0] Wgt_9_411, // sfix19_En18
  input [18:0] Wgt_9_412, // sfix19_En18
  input [18:0] Wgt_9_413, // sfix19_En18
  input [18:0] Wgt_9_414, // sfix19_En18
  input [18:0] Wgt_9_415, // sfix19_En18
  input [18:0] Wgt_9_416, // sfix19_En18
  input [18:0] Wgt_9_417, // sfix19_En18
  input [18:0] Wgt_9_418, // sfix19_En18
  input [18:0] Wgt_9_419, // sfix19_En18
  input [18:0] Wgt_9_420, // sfix19_En18
  input [18:0] Wgt_9_421, // sfix19_En18
  input [18:0] Wgt_9_422, // sfix19_En18
  input [18:0] Wgt_9_423, // sfix19_En18
  input [18:0] Wgt_9_424, // sfix19_En18
  input [18:0] Wgt_9_425, // sfix19_En18
  input [18:0] Wgt_9_426, // sfix19_En18
  input [18:0] Wgt_9_427, // sfix19_En18
  input [18:0] Wgt_9_428, // sfix19_En18
  input [18:0] Wgt_9_429, // sfix19_En18
  input [18:0] Wgt_9_430, // sfix19_En18
  input [18:0] Wgt_9_431, // sfix19_En18
  input [18:0] Wgt_9_432, // sfix19_En18
  input [18:0] Wgt_9_433, // sfix19_En18
  input [18:0] Wgt_9_434, // sfix19_En18
  input [18:0] Wgt_9_435, // sfix19_En18
  input [18:0] Wgt_9_436, // sfix19_En18
  input [18:0] Wgt_9_437, // sfix19_En18
  input [18:0] Wgt_9_438, // sfix19_En18
  input [18:0] Wgt_9_439, // sfix19_En18
  input [18:0] Wgt_9_440, // sfix19_En18
  input [18:0] Wgt_9_441, // sfix19_En18
  input [18:0] Wgt_9_442, // sfix19_En18
  input [18:0] Wgt_9_443, // sfix19_En18
  input [18:0] Wgt_9_444, // sfix19_En18
  input [18:0] Wgt_9_445, // sfix19_En18
  input [18:0] Wgt_9_446, // sfix19_En18
  input [18:0] Wgt_9_447, // sfix19_En18
  input [18:0] Wgt_9_448, // sfix19_En18
  input [18:0] Wgt_9_449, // sfix19_En18
  input [18:0] Wgt_9_450, // sfix19_En18
  input [18:0] Wgt_9_451, // sfix19_En18
  input [18:0] Wgt_9_452, // sfix19_En18
  input [18:0] Wgt_9_453, // sfix19_En18
  input [18:0] Wgt_9_454, // sfix19_En18
  input [18:0] Wgt_9_455, // sfix19_En18
  input [18:0] Wgt_9_456, // sfix19_En18
  input [18:0] Wgt_9_457, // sfix19_En18
  input [18:0] Wgt_9_458, // sfix19_En18
  input [18:0] Wgt_9_459, // sfix19_En18
  input [18:0] Wgt_9_460, // sfix19_En18
  input [18:0] Wgt_9_461, // sfix19_En18
  input [18:0] Wgt_9_462, // sfix19_En18
  input [18:0] Wgt_9_463, // sfix19_En18
  input [18:0] Wgt_9_464, // sfix19_En18
  input [18:0] Wgt_9_465, // sfix19_En18
  input [18:0] Wgt_9_466, // sfix19_En18
  input [18:0] Wgt_9_467, // sfix19_En18
  input [18:0] Wgt_9_468, // sfix19_En18
  input [18:0] Wgt_9_469, // sfix19_En18
  input [18:0] Wgt_9_470, // sfix19_En18
  input [18:0] Wgt_9_471, // sfix19_En18
  input [18:0] Wgt_9_472, // sfix19_En18
  input [18:0] Wgt_9_473, // sfix19_En18
  input [18:0] Wgt_9_474, // sfix19_En18
  input [18:0] Wgt_9_475, // sfix19_En18
  input [18:0] Wgt_9_476, // sfix19_En18
  input [18:0] Wgt_9_477, // sfix19_En18
  input [18:0] Wgt_9_478, // sfix19_En18
  input [18:0] Wgt_9_479, // sfix19_En18
  input [18:0] Wgt_9_480, // sfix19_En18
  input [18:0] Wgt_9_481, // sfix19_En18
  input [18:0] Wgt_9_482, // sfix19_En18
  input [18:0] Wgt_9_483, // sfix19_En18
  input [18:0] Wgt_9_484, // sfix19_En18
  input [18:0] Wgt_9_485, // sfix19_En18
  input [18:0] Wgt_9_486, // sfix19_En18
  input [18:0] Wgt_9_487, // sfix19_En18
  input [18:0] Wgt_9_488, // sfix19_En18
  input [18:0] Wgt_9_489, // sfix19_En18
  input [18:0] Wgt_9_490, // sfix19_En18
  input [18:0] Wgt_9_491, // sfix19_En18
  input [18:0] Wgt_9_492, // sfix19_En18
  input [18:0] Wgt_9_493, // sfix19_En18
  input [18:0] Wgt_9_494, // sfix19_En18
  input [18:0] Wgt_9_495, // sfix19_En18
  input [18:0] Wgt_9_496, // sfix19_En18
  input [18:0] Wgt_9_497, // sfix19_En18
  input [18:0] Wgt_9_498, // sfix19_En18
  input [18:0] Wgt_9_499, // sfix19_En18
  input [18:0] Wgt_9_500, // sfix19_En18
  input [18:0] Wgt_9_501, // sfix19_En18
  input [18:0] Wgt_9_502, // sfix19_En18
  input [18:0] Wgt_9_503, // sfix19_En18
  input [18:0] Wgt_9_504, // sfix19_En18
  input [18:0] Wgt_9_505, // sfix19_En18
  input [18:0] Wgt_9_506, // sfix19_En18
  input [18:0] Wgt_9_507, // sfix19_En18
  input [18:0] Wgt_9_508, // sfix19_En18
  input [18:0] Wgt_9_509, // sfix19_En18
  input [18:0] Wgt_9_510, // sfix19_En18
  input [18:0] Wgt_9_511, // sfix19_En18
  input [18:0] Wgt_9_512, // sfix19_En18
  input [18:0] Wgt_9_513, // sfix19_En18
  input [18:0] Wgt_9_514, // sfix19_En18
  input [18:0] Wgt_9_515, // sfix19_En18
  input [18:0] Wgt_9_516, // sfix19_En18
  input [18:0] Wgt_9_517, // sfix19_En18
  input [18:0] Wgt_9_518, // sfix19_En18
  input [18:0] Wgt_9_519, // sfix19_En18
  input [18:0] Wgt_9_520, // sfix19_En18
  input [18:0] Wgt_9_521, // sfix19_En18
  input [18:0] Wgt_9_522, // sfix19_En18
  input [18:0] Wgt_9_523, // sfix19_En18
  input [18:0] Wgt_9_524, // sfix19_En18
  input [18:0] Wgt_9_525, // sfix19_En18
  input [18:0] Wgt_9_526, // sfix19_En18
  input [18:0] Wgt_9_527, // sfix19_En18
  input [18:0] Wgt_9_528, // sfix19_En18
  input [18:0] Wgt_9_529, // sfix19_En18
  input [18:0] Wgt_9_530, // sfix19_En18
  input [18:0] Wgt_9_531, // sfix19_En18
  input [18:0] Wgt_9_532, // sfix19_En18
  input [18:0] Wgt_9_533, // sfix19_En18
  input [18:0] Wgt_9_534, // sfix19_En18
  input [18:0] Wgt_9_535, // sfix19_En18
  input [18:0] Wgt_9_536, // sfix19_En18
  input [18:0] Wgt_9_537, // sfix19_En18
  input [18:0] Wgt_9_538, // sfix19_En18
  input [18:0] Wgt_9_539, // sfix19_En18
  input [18:0] Wgt_9_540, // sfix19_En18
  input [18:0] Wgt_9_541, // sfix19_En18
  input [18:0] Wgt_9_542, // sfix19_En18
  input [18:0] Wgt_9_543, // sfix19_En18
  input [18:0] Wgt_9_544, // sfix19_En18
  input [18:0] Wgt_9_545, // sfix19_En18
  input [18:0] Wgt_9_546, // sfix19_En18
  input [18:0] Wgt_9_547, // sfix19_En18
  input [18:0] Wgt_9_548, // sfix19_En18
  input [18:0] Wgt_9_549, // sfix19_En18
  input [18:0] Wgt_9_550, // sfix19_En18
  input [18:0] Wgt_9_551, // sfix19_En18
  input [18:0] Wgt_9_552, // sfix19_En18
  input [18:0] Wgt_9_553, // sfix19_En18
  input [18:0] Wgt_9_554, // sfix19_En18
  input [18:0] Wgt_9_555, // sfix19_En18
  input [18:0] Wgt_9_556, // sfix19_En18
  input [18:0] Wgt_9_557, // sfix19_En18
  input [18:0] Wgt_9_558, // sfix19_En18
  input [18:0] Wgt_9_559, // sfix19_En18
  input [18:0] Wgt_9_560, // sfix19_En18
  input [18:0] Wgt_9_561, // sfix19_En18
  input [18:0] Wgt_9_562, // sfix19_En18
  input [18:0] Wgt_9_563, // sfix19_En18
  input [18:0] Wgt_9_564, // sfix19_En18
  input [18:0] Wgt_9_565, // sfix19_En18
  input [18:0] Wgt_9_566, // sfix19_En18
  input [18:0] Wgt_9_567, // sfix19_En18
  input [18:0] Wgt_9_568, // sfix19_En18
  input [18:0] Wgt_9_569, // sfix19_En18
  input [18:0] Wgt_9_570, // sfix19_En18
  input [18:0] Wgt_9_571, // sfix19_En18
  input [18:0] Wgt_9_572, // sfix19_En18
  input [18:0] Wgt_9_573, // sfix19_En18
  input [18:0] Wgt_9_574, // sfix19_En18
  input [18:0] Wgt_9_575, // sfix19_En18
  input [18:0] Wgt_9_576, // sfix19_En18
  input [18:0] Wgt_9_577, // sfix19_En18
  input [18:0] Wgt_9_578, // sfix19_En18
  input [18:0] Wgt_9_579, // sfix19_En18
  input [18:0] Wgt_9_580, // sfix19_En18
  input [18:0] Wgt_9_581, // sfix19_En18
  input [18:0] Wgt_9_582, // sfix19_En18
  input [18:0] Wgt_9_583, // sfix19_En18
  input [18:0] Wgt_9_584, // sfix19_En18
  input [18:0] Wgt_9_585, // sfix19_En18
  input [18:0] Wgt_9_586, // sfix19_En18
  input [18:0] Wgt_9_587, // sfix19_En18
  input [18:0] Wgt_9_588, // sfix19_En18
  input [18:0] Wgt_9_589, // sfix19_En18
  input [18:0] Wgt_9_590, // sfix19_En18
  input [18:0] Wgt_9_591, // sfix19_En18
  input [18:0] Wgt_9_592, // sfix19_En18
  input [18:0] Wgt_9_593, // sfix19_En18
  input [18:0] Wgt_9_594, // sfix19_En18
  input [18:0] Wgt_9_595, // sfix19_En18
  input [18:0] Wgt_9_596, // sfix19_En18
  input [18:0] Wgt_9_597, // sfix19_En18
  input [18:0] Wgt_9_598, // sfix19_En18
  input [18:0] Wgt_9_599, // sfix19_En18
  input [18:0] Wgt_9_600, // sfix19_En18
  input [18:0] Wgt_9_601, // sfix19_En18
  input [18:0] Wgt_9_602, // sfix19_En18
  input [18:0] Wgt_9_603, // sfix19_En18
  input [18:0] Wgt_9_604, // sfix19_En18
  input [18:0] Wgt_9_605, // sfix19_En18
  input [18:0] Wgt_9_606, // sfix19_En18
  input [18:0] Wgt_9_607, // sfix19_En18
  input [18:0] Wgt_9_608, // sfix19_En18
  input [18:0] Wgt_9_609, // sfix19_En18
  input [18:0] Wgt_9_610, // sfix19_En18
  input [18:0] Wgt_9_611, // sfix19_En18
  input [18:0] Wgt_9_612, // sfix19_En18
  input [18:0] Wgt_9_613, // sfix19_En18
  input [18:0] Wgt_9_614, // sfix19_En18
  input [18:0] Wgt_9_615, // sfix19_En18
  input [18:0] Wgt_9_616, // sfix19_En18
  input [18:0] Wgt_9_617, // sfix19_En18
  input [18:0] Wgt_9_618, // sfix19_En18
  input [18:0] Wgt_9_619, // sfix19_En18
  input [18:0] Wgt_9_620, // sfix19_En18
  input [18:0] Wgt_9_621, // sfix19_En18
  input [18:0] Wgt_9_622, // sfix19_En18
  input [18:0] Wgt_9_623, // sfix19_En18
  input [18:0] Wgt_9_624, // sfix19_En18
  input [18:0] Wgt_9_625, // sfix19_En18
  input [18:0] Wgt_9_626, // sfix19_En18
  input [18:0] Wgt_9_627, // sfix19_En18
  input [18:0] Wgt_9_628, // sfix19_En18
  input [18:0] Wgt_9_629, // sfix19_En18
  input [18:0] Wgt_9_630, // sfix19_En18
  input [18:0] Wgt_9_631, // sfix19_En18
  input [18:0] Wgt_9_632, // sfix19_En18
  input [18:0] Wgt_9_633, // sfix19_En18
  input [18:0] Wgt_9_634, // sfix19_En18
  input [18:0] Wgt_9_635, // sfix19_En18
  input [18:0] Wgt_9_636, // sfix19_En18
  input [18:0] Wgt_9_637, // sfix19_En18
  input [18:0] Wgt_9_638, // sfix19_En18
  input [18:0] Wgt_9_639, // sfix19_En18
  input [18:0] Wgt_9_640, // sfix19_En18
  input [18:0] Wgt_9_641, // sfix19_En18
  input [18:0] Wgt_9_642, // sfix19_En18
  input [18:0] Wgt_9_643, // sfix19_En18
  input [18:0] Wgt_9_644, // sfix19_En18
  input [18:0] Wgt_9_645, // sfix19_En18
  input [18:0] Wgt_9_646, // sfix19_En18
  input [18:0] Wgt_9_647, // sfix19_En18
  input [18:0] Wgt_9_648, // sfix19_En18
  input [18:0] Wgt_9_649, // sfix19_En18
  input [18:0] Wgt_9_650, // sfix19_En18
  input [18:0] Wgt_9_651, // sfix19_En18
  input [18:0] Wgt_9_652, // sfix19_En18
  input [18:0] Wgt_9_653, // sfix19_En18
  input [18:0] Wgt_9_654, // sfix19_En18
  input [18:0] Wgt_9_655, // sfix19_En18
  input [18:0] Wgt_9_656, // sfix19_En18
  input [18:0] Wgt_9_657, // sfix19_En18
  input [18:0] Wgt_9_658, // sfix19_En18
  input [18:0] Wgt_9_659, // sfix19_En18
  input [18:0] Wgt_9_660, // sfix19_En18
  input [18:0] Wgt_9_661, // sfix19_En18
  input [18:0] Wgt_9_662, // sfix19_En18
  input [18:0] Wgt_9_663, // sfix19_En18
  input [18:0] Wgt_9_664, // sfix19_En18
  input [18:0] Wgt_9_665, // sfix19_En18
  input [18:0] Wgt_9_666, // sfix19_En18
  input [18:0] Wgt_9_667, // sfix19_En18
  input [18:0] Wgt_9_668, // sfix19_En18
  input [18:0] Wgt_9_669, // sfix19_En18
  input [18:0] Wgt_9_670, // sfix19_En18
  input [18:0] Wgt_9_671, // sfix19_En18
  input [18:0] Wgt_9_672, // sfix19_En18
  input [18:0] Wgt_9_673, // sfix19_En18
  input [18:0] Wgt_9_674, // sfix19_En18
  input [18:0] Wgt_9_675, // sfix19_En18
  input [18:0] Wgt_9_676, // sfix19_En18
  input [18:0] Wgt_9_677, // sfix19_En18
  input [18:0] Wgt_9_678, // sfix19_En18
  input [18:0] Wgt_9_679, // sfix19_En18
  input [18:0] Wgt_9_680, // sfix19_En18
  input [18:0] Wgt_9_681, // sfix19_En18
  input [18:0] Wgt_9_682, // sfix19_En18
  input [18:0] Wgt_9_683, // sfix19_En18
  input [18:0] Wgt_9_684, // sfix19_En18
  input [18:0] Wgt_9_685, // sfix19_En18
  input [18:0] Wgt_9_686, // sfix19_En18
  input [18:0] Wgt_9_687, // sfix19_En18
  input [18:0] Wgt_9_688, // sfix19_En18
  input [18:0] Wgt_9_689, // sfix19_En18
  input [18:0] Wgt_9_690, // sfix19_En18
  input [18:0] Wgt_9_691, // sfix19_En18
  input [18:0] Wgt_9_692, // sfix19_En18
  input [18:0] Wgt_9_693, // sfix19_En18
  input [18:0] Wgt_9_694, // sfix19_En18
  input [18:0] Wgt_9_695, // sfix19_En18
  input [18:0] Wgt_9_696, // sfix19_En18
  input [18:0] Wgt_9_697, // sfix19_En18
  input [18:0] Wgt_9_698, // sfix19_En18
  input [18:0] Wgt_9_699, // sfix19_En18
  input [18:0] Wgt_9_700, // sfix19_En18
  input [18:0] Wgt_9_701, // sfix19_En18
  input [18:0] Wgt_9_702, // sfix19_En18
  input [18:0] Wgt_9_703, // sfix19_En18
  input [18:0] Wgt_9_704, // sfix19_En18
  input [18:0] Wgt_9_705, // sfix19_En18
  input [18:0] Wgt_9_706, // sfix19_En18
  input [18:0] Wgt_9_707, // sfix19_En18
  input [18:0] Wgt_9_708, // sfix19_En18
  input [18:0] Wgt_9_709, // sfix19_En18
  input [18:0] Wgt_9_710, // sfix19_En18
  input [18:0] Wgt_9_711, // sfix19_En18
  input [18:0] Wgt_9_712, // sfix19_En18
  input [18:0] Wgt_9_713, // sfix19_En18
  input [18:0] Wgt_9_714, // sfix19_En18
  input [18:0] Wgt_9_715, // sfix19_En18
  input [18:0] Wgt_9_716, // sfix19_En18
  input [18:0] Wgt_9_717, // sfix19_En18
  input [18:0] Wgt_9_718, // sfix19_En18
  input [18:0] Wgt_9_719, // sfix19_En18
  input [18:0] Wgt_9_720, // sfix19_En18
  input [18:0] Wgt_9_721, // sfix19_En18
  input [18:0] Wgt_9_722, // sfix19_En18
  input [18:0] Wgt_9_723, // sfix19_En18
  input [18:0] Wgt_9_724, // sfix19_En18
  input [18:0] Wgt_9_725, // sfix19_En18
  input [18:0] Wgt_9_726, // sfix19_En18
  input [18:0] Wgt_9_727, // sfix19_En18
  input [18:0] Wgt_9_728, // sfix19_En18
  input [18:0] Wgt_9_729, // sfix19_En18
  input [18:0] Wgt_9_730, // sfix19_En18
  input [18:0] Wgt_9_731, // sfix19_En18
  input [18:0] Wgt_9_732, // sfix19_En18
  input [18:0] Wgt_9_733, // sfix19_En18
  input [18:0] Wgt_9_734, // sfix19_En18
  input [18:0] Wgt_9_735, // sfix19_En18
  input [18:0] Wgt_9_736, // sfix19_En18
  input [18:0] Wgt_9_737, // sfix19_En18
  input [18:0] Wgt_9_738, // sfix19_En18
  input [18:0] Wgt_9_739, // sfix19_En18
  input [18:0] Wgt_9_740, // sfix19_En18
  input [18:0] Wgt_9_741, // sfix19_En18
  input [18:0] Wgt_9_742, // sfix19_En18
  input [18:0] Wgt_9_743, // sfix19_En18
  input [18:0] Wgt_9_744, // sfix19_En18
  input [18:0] Wgt_9_745, // sfix19_En18
  input [18:0] Wgt_9_746, // sfix19_En18
  input [18:0] Wgt_9_747, // sfix19_En18
  input [18:0] Wgt_9_748, // sfix19_En18
  input [18:0] Wgt_9_749, // sfix19_En18
  input [18:0] Wgt_9_750, // sfix19_En18
  input [18:0] Wgt_9_751, // sfix19_En18
  input [18:0] Wgt_9_752, // sfix19_En18
  input [18:0] Wgt_9_753, // sfix19_En18
  input [18:0] Wgt_9_754, // sfix19_En18
  input [18:0] Wgt_9_755, // sfix19_En18
  input [18:0] Wgt_9_756, // sfix19_En18
  input [18:0] Wgt_9_757, // sfix19_En18
  input [18:0] Wgt_9_758, // sfix19_En18
  input [18:0] Wgt_9_759, // sfix19_En18
  input [18:0] Wgt_9_760, // sfix19_En18
  input [18:0] Wgt_9_761, // sfix19_En18
  input [18:0] Wgt_9_762, // sfix19_En18
  input [18:0] Wgt_9_763, // sfix19_En18
  input [18:0] Wgt_9_764, // sfix19_En18
  input [18:0] Wgt_9_765, // sfix19_En18
  input [18:0] Wgt_9_766, // sfix19_En18
  input [18:0] Wgt_9_767, // sfix19_En18
  input [18:0] Wgt_9_768, // sfix19_En18
  input [18:0] Wgt_9_769, // sfix19_En18
  input [18:0] Wgt_9_770, // sfix19_En18
  input [18:0] Wgt_9_771, // sfix19_En18
  input [18:0] Wgt_9_772, // sfix19_En18
  input [18:0] Wgt_9_773, // sfix19_En18
  input [18:0] Wgt_9_774, // sfix19_En18
  input [18:0] Wgt_9_775, // sfix19_En18
  input [18:0] Wgt_9_776, // sfix19_En18
  input [18:0] Wgt_9_777, // sfix19_En18
  input [18:0] Wgt_9_778, // sfix19_En18
  input [18:0] Wgt_9_779, // sfix19_En18
  input [18:0] Wgt_9_780, // sfix19_En18
  input [18:0] Wgt_9_781, // sfix19_En18
  input [18:0] Wgt_9_782, // sfix19_En18
  input [18:0] Wgt_9_783, // sfix19_En18
  input [18:0] Wgt_9_784, // sfix19_En18
 input [9:0] Pix_0, // sfix10_En0
 input [9:0] Pix_1, // sfix10_En0
 input [9:0] Pix_2, // sfix10_En0
 input [9:0] Pix_3, // sfix10_En0
 input [9:0] Pix_4, // sfix10_En0
 input [9:0] Pix_5, // sfix10_En0
 input [9:0] Pix_6, // sfix10_En0
 input [9:0] Pix_7, // sfix10_En0
 input [9:0] Pix_8, // sfix10_En0
 input [9:0] Pix_9, // sfix10_En0
 input [9:0] Pix_10, // sfix10_En0
 input [9:0] Pix_11, // sfix10_En0
 input [9:0] Pix_12, // sfix10_En0
 input [9:0] Pix_13, // sfix10_En0
 input [9:0] Pix_14, // sfix10_En0
 input [9:0] Pix_15, // sfix10_En0
 input [9:0] Pix_16, // sfix10_En0
 input [9:0] Pix_17, // sfix10_En0
 input [9:0] Pix_18, // sfix10_En0
 input [9:0] Pix_19, // sfix10_En0
 input [9:0] Pix_20, // sfix10_En0
 input [9:0] Pix_21, // sfix10_En0
 input [9:0] Pix_22, // sfix10_En0
 input [9:0] Pix_23, // sfix10_En0
 input [9:0] Pix_24, // sfix10_En0
 input [9:0] Pix_25, // sfix10_En0
 input [9:0] Pix_26, // sfix10_En0
 input [9:0] Pix_27, // sfix10_En0
 input [9:0] Pix_28, // sfix10_En0
 input [9:0] Pix_29, // sfix10_En0
 input [9:0] Pix_30, // sfix10_En0
 input [9:0] Pix_31, // sfix10_En0
 input [9:0] Pix_32, // sfix10_En0
 input [9:0] Pix_33, // sfix10_En0
 input [9:0] Pix_34, // sfix10_En0
 input [9:0] Pix_35, // sfix10_En0
 input [9:0] Pix_36, // sfix10_En0
 input [9:0] Pix_37, // sfix10_En0
 input [9:0] Pix_38, // sfix10_En0
 input [9:0] Pix_39, // sfix10_En0
 input [9:0] Pix_40, // sfix10_En0
 input [9:0] Pix_41, // sfix10_En0
 input [9:0] Pix_42, // sfix10_En0
 input [9:0] Pix_43, // sfix10_En0
 input [9:0] Pix_44, // sfix10_En0
 input [9:0] Pix_45, // sfix10_En0
 input [9:0] Pix_46, // sfix10_En0
 input [9:0] Pix_47, // sfix10_En0
 input [9:0] Pix_48, // sfix10_En0
 input [9:0] Pix_49, // sfix10_En0
 input [9:0] Pix_50, // sfix10_En0
 input [9:0] Pix_51, // sfix10_En0
 input [9:0] Pix_52, // sfix10_En0
 input [9:0] Pix_53, // sfix10_En0
 input [9:0] Pix_54, // sfix10_En0
 input [9:0] Pix_55, // sfix10_En0
 input [9:0] Pix_56, // sfix10_En0
 input [9:0] Pix_57, // sfix10_En0
 input [9:0] Pix_58, // sfix10_En0
 input [9:0] Pix_59, // sfix10_En0
 input [9:0] Pix_60, // sfix10_En0
 input [9:0] Pix_61, // sfix10_En0
 input [9:0] Pix_62, // sfix10_En0
 input [9:0] Pix_63, // sfix10_En0
 input [9:0] Pix_64, // sfix10_En0
 input [9:0] Pix_65, // sfix10_En0
 input [9:0] Pix_66, // sfix10_En0
 input [9:0] Pix_67, // sfix10_En0
 input [9:0] Pix_68, // sfix10_En0
 input [9:0] Pix_69, // sfix10_En0
 input [9:0] Pix_70, // sfix10_En0
 input [9:0] Pix_71, // sfix10_En0
 input [9:0] Pix_72, // sfix10_En0
 input [9:0] Pix_73, // sfix10_En0
 input [9:0] Pix_74, // sfix10_En0
 input [9:0] Pix_75, // sfix10_En0
 input [9:0] Pix_76, // sfix10_En0
 input [9:0] Pix_77, // sfix10_En0
 input [9:0] Pix_78, // sfix10_En0
 input [9:0] Pix_79, // sfix10_En0
 input [9:0] Pix_80, // sfix10_En0
 input [9:0] Pix_81, // sfix10_En0
 input [9:0] Pix_82, // sfix10_En0
 input [9:0] Pix_83, // sfix10_En0
 input [9:0] Pix_84, // sfix10_En0
 input [9:0] Pix_85, // sfix10_En0
 input [9:0] Pix_86, // sfix10_En0
 input [9:0] Pix_87, // sfix10_En0
 input [9:0] Pix_88, // sfix10_En0
 input [9:0] Pix_89, // sfix10_En0
 input [9:0] Pix_90, // sfix10_En0
 input [9:0] Pix_91, // sfix10_En0
 input [9:0] Pix_92, // sfix10_En0
 input [9:0] Pix_93, // sfix10_En0
 input [9:0] Pix_94, // sfix10_En0
 input [9:0] Pix_95, // sfix10_En0
 input [9:0] Pix_96, // sfix10_En0
 input [9:0] Pix_97, // sfix10_En0
 input [9:0] Pix_98, // sfix10_En0
 input [9:0] Pix_99, // sfix10_En0
 input [9:0] Pix_100, // sfix10_En0
 input [9:0] Pix_101, // sfix10_En0
 input [9:0] Pix_102, // sfix10_En0
 input [9:0] Pix_103, // sfix10_En0
 input [9:0] Pix_104, // sfix10_En0
 input [9:0] Pix_105, // sfix10_En0
 input [9:0] Pix_106, // sfix10_En0
 input [9:0] Pix_107, // sfix10_En0
 input [9:0] Pix_108, // sfix10_En0
 input [9:0] Pix_109, // sfix10_En0
 input [9:0] Pix_110, // sfix10_En0
 input [9:0] Pix_111, // sfix10_En0
 input [9:0] Pix_112, // sfix10_En0
 input [9:0] Pix_113, // sfix10_En0
 input [9:0] Pix_114, // sfix10_En0
 input [9:0] Pix_115, // sfix10_En0
 input [9:0] Pix_116, // sfix10_En0
 input [9:0] Pix_117, // sfix10_En0
 input [9:0] Pix_118, // sfix10_En0
 input [9:0] Pix_119, // sfix10_En0
 input [9:0] Pix_120, // sfix10_En0
 input [9:0] Pix_121, // sfix10_En0
 input [9:0] Pix_122, // sfix10_En0
 input [9:0] Pix_123, // sfix10_En0
 input [9:0] Pix_124, // sfix10_En0
 input [9:0] Pix_125, // sfix10_En0
 input [9:0] Pix_126, // sfix10_En0
 input [9:0] Pix_127, // sfix10_En0
 input [9:0] Pix_128, // sfix10_En0
 input [9:0] Pix_129, // sfix10_En0
 input [9:0] Pix_130, // sfix10_En0
 input [9:0] Pix_131, // sfix10_En0
 input [9:0] Pix_132, // sfix10_En0
 input [9:0] Pix_133, // sfix10_En0
 input [9:0] Pix_134, // sfix10_En0
 input [9:0] Pix_135, // sfix10_En0
 input [9:0] Pix_136, // sfix10_En0
 input [9:0] Pix_137, // sfix10_En0
 input [9:0] Pix_138, // sfix10_En0
 input [9:0] Pix_139, // sfix10_En0
 input [9:0] Pix_140, // sfix10_En0
 input [9:0] Pix_141, // sfix10_En0
 input [9:0] Pix_142, // sfix10_En0
 input [9:0] Pix_143, // sfix10_En0
 input [9:0] Pix_144, // sfix10_En0
 input [9:0] Pix_145, // sfix10_En0
 input [9:0] Pix_146, // sfix10_En0
 input [9:0] Pix_147, // sfix10_En0
 input [9:0] Pix_148, // sfix10_En0
 input [9:0] Pix_149, // sfix10_En0
 input [9:0] Pix_150, // sfix10_En0
 input [9:0] Pix_151, // sfix10_En0
 input [9:0] Pix_152, // sfix10_En0
 input [9:0] Pix_153, // sfix10_En0
 input [9:0] Pix_154, // sfix10_En0
 input [9:0] Pix_155, // sfix10_En0
 input [9:0] Pix_156, // sfix10_En0
 input [9:0] Pix_157, // sfix10_En0
 input [9:0] Pix_158, // sfix10_En0
 input [9:0] Pix_159, // sfix10_En0
 input [9:0] Pix_160, // sfix10_En0
 input [9:0] Pix_161, // sfix10_En0
 input [9:0] Pix_162, // sfix10_En0
 input [9:0] Pix_163, // sfix10_En0
 input [9:0] Pix_164, // sfix10_En0
 input [9:0] Pix_165, // sfix10_En0
 input [9:0] Pix_166, // sfix10_En0
 input [9:0] Pix_167, // sfix10_En0
 input [9:0] Pix_168, // sfix10_En0
 input [9:0] Pix_169, // sfix10_En0
 input [9:0] Pix_170, // sfix10_En0
 input [9:0] Pix_171, // sfix10_En0
 input [9:0] Pix_172, // sfix10_En0
 input [9:0] Pix_173, // sfix10_En0
 input [9:0] Pix_174, // sfix10_En0
 input [9:0] Pix_175, // sfix10_En0
 input [9:0] Pix_176, // sfix10_En0
 input [9:0] Pix_177, // sfix10_En0
 input [9:0] Pix_178, // sfix10_En0
 input [9:0] Pix_179, // sfix10_En0
 input [9:0] Pix_180, // sfix10_En0
 input [9:0] Pix_181, // sfix10_En0
 input [9:0] Pix_182, // sfix10_En0
 input [9:0] Pix_183, // sfix10_En0
 input [9:0] Pix_184, // sfix10_En0
 input [9:0] Pix_185, // sfix10_En0
 input [9:0] Pix_186, // sfix10_En0
 input [9:0] Pix_187, // sfix10_En0
 input [9:0] Pix_188, // sfix10_En0
 input [9:0] Pix_189, // sfix10_En0
 input [9:0] Pix_190, // sfix10_En0
 input [9:0] Pix_191, // sfix10_En0
 input [9:0] Pix_192, // sfix10_En0
 input [9:0] Pix_193, // sfix10_En0
 input [9:0] Pix_194, // sfix10_En0
 input [9:0] Pix_195, // sfix10_En0
 input [9:0] Pix_196, // sfix10_En0
 input [9:0] Pix_197, // sfix10_En0
 input [9:0] Pix_198, // sfix10_En0
 input [9:0] Pix_199, // sfix10_En0
 input [9:0] Pix_200, // sfix10_En0
 input [9:0] Pix_201, // sfix10_En0
 input [9:0] Pix_202, // sfix10_En0
 input [9:0] Pix_203, // sfix10_En0
 input [9:0] Pix_204, // sfix10_En0
 input [9:0] Pix_205, // sfix10_En0
 input [9:0] Pix_206, // sfix10_En0
 input [9:0] Pix_207, // sfix10_En0
 input [9:0] Pix_208, // sfix10_En0
 input [9:0] Pix_209, // sfix10_En0
 input [9:0] Pix_210, // sfix10_En0
 input [9:0] Pix_211, // sfix10_En0
 input [9:0] Pix_212, // sfix10_En0
 input [9:0] Pix_213, // sfix10_En0
 input [9:0] Pix_214, // sfix10_En0
 input [9:0] Pix_215, // sfix10_En0
 input [9:0] Pix_216, // sfix10_En0
 input [9:0] Pix_217, // sfix10_En0
 input [9:0] Pix_218, // sfix10_En0
 input [9:0] Pix_219, // sfix10_En0
 input [9:0] Pix_220, // sfix10_En0
 input [9:0] Pix_221, // sfix10_En0
 input [9:0] Pix_222, // sfix10_En0
 input [9:0] Pix_223, // sfix10_En0
 input [9:0] Pix_224, // sfix10_En0
 input [9:0] Pix_225, // sfix10_En0
 input [9:0] Pix_226, // sfix10_En0
 input [9:0] Pix_227, // sfix10_En0
 input [9:0] Pix_228, // sfix10_En0
 input [9:0] Pix_229, // sfix10_En0
 input [9:0] Pix_230, // sfix10_En0
 input [9:0] Pix_231, // sfix10_En0
 input [9:0] Pix_232, // sfix10_En0
 input [9:0] Pix_233, // sfix10_En0
 input [9:0] Pix_234, // sfix10_En0
 input [9:0] Pix_235, // sfix10_En0
 input [9:0] Pix_236, // sfix10_En0
 input [9:0] Pix_237, // sfix10_En0
 input [9:0] Pix_238, // sfix10_En0
 input [9:0] Pix_239, // sfix10_En0
 input [9:0] Pix_240, // sfix10_En0
 input [9:0] Pix_241, // sfix10_En0
 input [9:0] Pix_242, // sfix10_En0
 input [9:0] Pix_243, // sfix10_En0
 input [9:0] Pix_244, // sfix10_En0
 input [9:0] Pix_245, // sfix10_En0
 input [9:0] Pix_246, // sfix10_En0
 input [9:0] Pix_247, // sfix10_En0
 input [9:0] Pix_248, // sfix10_En0
 input [9:0] Pix_249, // sfix10_En0
 input [9:0] Pix_250, // sfix10_En0
 input [9:0] Pix_251, // sfix10_En0
 input [9:0] Pix_252, // sfix10_En0
 input [9:0] Pix_253, // sfix10_En0
 input [9:0] Pix_254, // sfix10_En0
 input [9:0] Pix_255, // sfix10_En0
 input [9:0] Pix_256, // sfix10_En0
 input [9:0] Pix_257, // sfix10_En0
 input [9:0] Pix_258, // sfix10_En0
 input [9:0] Pix_259, // sfix10_En0
 input [9:0] Pix_260, // sfix10_En0
 input [9:0] Pix_261, // sfix10_En0
 input [9:0] Pix_262, // sfix10_En0
 input [9:0] Pix_263, // sfix10_En0
 input [9:0] Pix_264, // sfix10_En0
 input [9:0] Pix_265, // sfix10_En0
 input [9:0] Pix_266, // sfix10_En0
 input [9:0] Pix_267, // sfix10_En0
 input [9:0] Pix_268, // sfix10_En0
 input [9:0] Pix_269, // sfix10_En0
 input [9:0] Pix_270, // sfix10_En0
 input [9:0] Pix_271, // sfix10_En0
 input [9:0] Pix_272, // sfix10_En0
 input [9:0] Pix_273, // sfix10_En0
 input [9:0] Pix_274, // sfix10_En0
 input [9:0] Pix_275, // sfix10_En0
 input [9:0] Pix_276, // sfix10_En0
 input [9:0] Pix_277, // sfix10_En0
 input [9:0] Pix_278, // sfix10_En0
 input [9:0] Pix_279, // sfix10_En0
 input [9:0] Pix_280, // sfix10_En0
 input [9:0] Pix_281, // sfix10_En0
 input [9:0] Pix_282, // sfix10_En0
 input [9:0] Pix_283, // sfix10_En0
 input [9:0] Pix_284, // sfix10_En0
 input [9:0] Pix_285, // sfix10_En0
 input [9:0] Pix_286, // sfix10_En0
 input [9:0] Pix_287, // sfix10_En0
 input [9:0] Pix_288, // sfix10_En0
 input [9:0] Pix_289, // sfix10_En0
 input [9:0] Pix_290, // sfix10_En0
 input [9:0] Pix_291, // sfix10_En0
 input [9:0] Pix_292, // sfix10_En0
 input [9:0] Pix_293, // sfix10_En0
 input [9:0] Pix_294, // sfix10_En0
 input [9:0] Pix_295, // sfix10_En0
 input [9:0] Pix_296, // sfix10_En0
 input [9:0] Pix_297, // sfix10_En0
 input [9:0] Pix_298, // sfix10_En0
 input [9:0] Pix_299, // sfix10_En0
 input [9:0] Pix_300, // sfix10_En0
 input [9:0] Pix_301, // sfix10_En0
 input [9:0] Pix_302, // sfix10_En0
 input [9:0] Pix_303, // sfix10_En0
 input [9:0] Pix_304, // sfix10_En0
 input [9:0] Pix_305, // sfix10_En0
 input [9:0] Pix_306, // sfix10_En0
 input [9:0] Pix_307, // sfix10_En0
 input [9:0] Pix_308, // sfix10_En0
 input [9:0] Pix_309, // sfix10_En0
 input [9:0] Pix_310, // sfix10_En0
 input [9:0] Pix_311, // sfix10_En0
 input [9:0] Pix_312, // sfix10_En0
 input [9:0] Pix_313, // sfix10_En0
 input [9:0] Pix_314, // sfix10_En0
 input [9:0] Pix_315, // sfix10_En0
 input [9:0] Pix_316, // sfix10_En0
 input [9:0] Pix_317, // sfix10_En0
 input [9:0] Pix_318, // sfix10_En0
 input [9:0] Pix_319, // sfix10_En0
 input [9:0] Pix_320, // sfix10_En0
 input [9:0] Pix_321, // sfix10_En0
 input [9:0] Pix_322, // sfix10_En0
 input [9:0] Pix_323, // sfix10_En0
 input [9:0] Pix_324, // sfix10_En0
 input [9:0] Pix_325, // sfix10_En0
 input [9:0] Pix_326, // sfix10_En0
 input [9:0] Pix_327, // sfix10_En0
 input [9:0] Pix_328, // sfix10_En0
 input [9:0] Pix_329, // sfix10_En0
 input [9:0] Pix_330, // sfix10_En0
 input [9:0] Pix_331, // sfix10_En0
 input [9:0] Pix_332, // sfix10_En0
 input [9:0] Pix_333, // sfix10_En0
 input [9:0] Pix_334, // sfix10_En0
 input [9:0] Pix_335, // sfix10_En0
 input [9:0] Pix_336, // sfix10_En0
 input [9:0] Pix_337, // sfix10_En0
 input [9:0] Pix_338, // sfix10_En0
 input [9:0] Pix_339, // sfix10_En0
 input [9:0] Pix_340, // sfix10_En0
 input [9:0] Pix_341, // sfix10_En0
 input [9:0] Pix_342, // sfix10_En0
 input [9:0] Pix_343, // sfix10_En0
 input [9:0] Pix_344, // sfix10_En0
 input [9:0] Pix_345, // sfix10_En0
 input [9:0] Pix_346, // sfix10_En0
 input [9:0] Pix_347, // sfix10_En0
 input [9:0] Pix_348, // sfix10_En0
 input [9:0] Pix_349, // sfix10_En0
 input [9:0] Pix_350, // sfix10_En0
 input [9:0] Pix_351, // sfix10_En0
 input [9:0] Pix_352, // sfix10_En0
 input [9:0] Pix_353, // sfix10_En0
 input [9:0] Pix_354, // sfix10_En0
 input [9:0] Pix_355, // sfix10_En0
 input [9:0] Pix_356, // sfix10_En0
 input [9:0] Pix_357, // sfix10_En0
 input [9:0] Pix_358, // sfix10_En0
 input [9:0] Pix_359, // sfix10_En0
 input [9:0] Pix_360, // sfix10_En0
 input [9:0] Pix_361, // sfix10_En0
 input [9:0] Pix_362, // sfix10_En0
 input [9:0] Pix_363, // sfix10_En0
 input [9:0] Pix_364, // sfix10_En0
 input [9:0] Pix_365, // sfix10_En0
 input [9:0] Pix_366, // sfix10_En0
 input [9:0] Pix_367, // sfix10_En0
 input [9:0] Pix_368, // sfix10_En0
 input [9:0] Pix_369, // sfix10_En0
 input [9:0] Pix_370, // sfix10_En0
 input [9:0] Pix_371, // sfix10_En0
 input [9:0] Pix_372, // sfix10_En0
 input [9:0] Pix_373, // sfix10_En0
 input [9:0] Pix_374, // sfix10_En0
 input [9:0] Pix_375, // sfix10_En0
 input [9:0] Pix_376, // sfix10_En0
 input [9:0] Pix_377, // sfix10_En0
 input [9:0] Pix_378, // sfix10_En0
 input [9:0] Pix_379, // sfix10_En0
 input [9:0] Pix_380, // sfix10_En0
 input [9:0] Pix_381, // sfix10_En0
 input [9:0] Pix_382, // sfix10_En0
 input [9:0] Pix_383, // sfix10_En0
 input [9:0] Pix_384, // sfix10_En0
 input [9:0] Pix_385, // sfix10_En0
 input [9:0] Pix_386, // sfix10_En0
 input [9:0] Pix_387, // sfix10_En0
 input [9:0] Pix_388, // sfix10_En0
 input [9:0] Pix_389, // sfix10_En0
 input [9:0] Pix_390, // sfix10_En0
 input [9:0] Pix_391, // sfix10_En0
 input [9:0] Pix_392, // sfix10_En0
 input [9:0] Pix_393, // sfix10_En0
 input [9:0] Pix_394, // sfix10_En0
 input [9:0] Pix_395, // sfix10_En0
 input [9:0] Pix_396, // sfix10_En0
 input [9:0] Pix_397, // sfix10_En0
 input [9:0] Pix_398, // sfix10_En0
 input [9:0] Pix_399, // sfix10_En0
 input [9:0] Pix_400, // sfix10_En0
 input [9:0] Pix_401, // sfix10_En0
 input [9:0] Pix_402, // sfix10_En0
 input [9:0] Pix_403, // sfix10_En0
 input [9:0] Pix_404, // sfix10_En0
 input [9:0] Pix_405, // sfix10_En0
 input [9:0] Pix_406, // sfix10_En0
 input [9:0] Pix_407, // sfix10_En0
 input [9:0] Pix_408, // sfix10_En0
 input [9:0] Pix_409, // sfix10_En0
 input [9:0] Pix_410, // sfix10_En0
 input [9:0] Pix_411, // sfix10_En0
 input [9:0] Pix_412, // sfix10_En0
 input [9:0] Pix_413, // sfix10_En0
 input [9:0] Pix_414, // sfix10_En0
 input [9:0] Pix_415, // sfix10_En0
 input [9:0] Pix_416, // sfix10_En0
 input [9:0] Pix_417, // sfix10_En0
 input [9:0] Pix_418, // sfix10_En0
 input [9:0] Pix_419, // sfix10_En0
 input [9:0] Pix_420, // sfix10_En0
 input [9:0] Pix_421, // sfix10_En0
 input [9:0] Pix_422, // sfix10_En0
 input [9:0] Pix_423, // sfix10_En0
 input [9:0] Pix_424, // sfix10_En0
 input [9:0] Pix_425, // sfix10_En0
 input [9:0] Pix_426, // sfix10_En0
 input [9:0] Pix_427, // sfix10_En0
 input [9:0] Pix_428, // sfix10_En0
 input [9:0] Pix_429, // sfix10_En0
 input [9:0] Pix_430, // sfix10_En0
 input [9:0] Pix_431, // sfix10_En0
 input [9:0] Pix_432, // sfix10_En0
 input [9:0] Pix_433, // sfix10_En0
 input [9:0] Pix_434, // sfix10_En0
 input [9:0] Pix_435, // sfix10_En0
 input [9:0] Pix_436, // sfix10_En0
 input [9:0] Pix_437, // sfix10_En0
 input [9:0] Pix_438, // sfix10_En0
 input [9:0] Pix_439, // sfix10_En0
 input [9:0] Pix_440, // sfix10_En0
 input [9:0] Pix_441, // sfix10_En0
 input [9:0] Pix_442, // sfix10_En0
 input [9:0] Pix_443, // sfix10_En0
 input [9:0] Pix_444, // sfix10_En0
 input [9:0] Pix_445, // sfix10_En0
 input [9:0] Pix_446, // sfix10_En0
 input [9:0] Pix_447, // sfix10_En0
 input [9:0] Pix_448, // sfix10_En0
 input [9:0] Pix_449, // sfix10_En0
 input [9:0] Pix_450, // sfix10_En0
 input [9:0] Pix_451, // sfix10_En0
 input [9:0] Pix_452, // sfix10_En0
 input [9:0] Pix_453, // sfix10_En0
 input [9:0] Pix_454, // sfix10_En0
 input [9:0] Pix_455, // sfix10_En0
 input [9:0] Pix_456, // sfix10_En0
 input [9:0] Pix_457, // sfix10_En0
 input [9:0] Pix_458, // sfix10_En0
 input [9:0] Pix_459, // sfix10_En0
 input [9:0] Pix_460, // sfix10_En0
 input [9:0] Pix_461, // sfix10_En0
 input [9:0] Pix_462, // sfix10_En0
 input [9:0] Pix_463, // sfix10_En0
 input [9:0] Pix_464, // sfix10_En0
 input [9:0] Pix_465, // sfix10_En0
 input [9:0] Pix_466, // sfix10_En0
 input [9:0] Pix_467, // sfix10_En0
 input [9:0] Pix_468, // sfix10_En0
 input [9:0] Pix_469, // sfix10_En0
 input [9:0] Pix_470, // sfix10_En0
 input [9:0] Pix_471, // sfix10_En0
 input [9:0] Pix_472, // sfix10_En0
 input [9:0] Pix_473, // sfix10_En0
 input [9:0] Pix_474, // sfix10_En0
 input [9:0] Pix_475, // sfix10_En0
 input [9:0] Pix_476, // sfix10_En0
 input [9:0] Pix_477, // sfix10_En0
 input [9:0] Pix_478, // sfix10_En0
 input [9:0] Pix_479, // sfix10_En0
 input [9:0] Pix_480, // sfix10_En0
 input [9:0] Pix_481, // sfix10_En0
 input [9:0] Pix_482, // sfix10_En0
 input [9:0] Pix_483, // sfix10_En0
 input [9:0] Pix_484, // sfix10_En0
 input [9:0] Pix_485, // sfix10_En0
 input [9:0] Pix_486, // sfix10_En0
 input [9:0] Pix_487, // sfix10_En0
 input [9:0] Pix_488, // sfix10_En0
 input [9:0] Pix_489, // sfix10_En0
 input [9:0] Pix_490, // sfix10_En0
 input [9:0] Pix_491, // sfix10_En0
 input [9:0] Pix_492, // sfix10_En0
 input [9:0] Pix_493, // sfix10_En0
 input [9:0] Pix_494, // sfix10_En0
 input [9:0] Pix_495, // sfix10_En0
 input [9:0] Pix_496, // sfix10_En0
 input [9:0] Pix_497, // sfix10_En0
 input [9:0] Pix_498, // sfix10_En0
 input [9:0] Pix_499, // sfix10_En0
 input [9:0] Pix_500, // sfix10_En0
 input [9:0] Pix_501, // sfix10_En0
 input [9:0] Pix_502, // sfix10_En0
 input [9:0] Pix_503, // sfix10_En0
 input [9:0] Pix_504, // sfix10_En0
 input [9:0] Pix_505, // sfix10_En0
 input [9:0] Pix_506, // sfix10_En0
 input [9:0] Pix_507, // sfix10_En0
 input [9:0] Pix_508, // sfix10_En0
 input [9:0] Pix_509, // sfix10_En0
 input [9:0] Pix_510, // sfix10_En0
 input [9:0] Pix_511, // sfix10_En0
 input [9:0] Pix_512, // sfix10_En0
 input [9:0] Pix_513, // sfix10_En0
 input [9:0] Pix_514, // sfix10_En0
 input [9:0] Pix_515, // sfix10_En0
 input [9:0] Pix_516, // sfix10_En0
 input [9:0] Pix_517, // sfix10_En0
 input [9:0] Pix_518, // sfix10_En0
 input [9:0] Pix_519, // sfix10_En0
 input [9:0] Pix_520, // sfix10_En0
 input [9:0] Pix_521, // sfix10_En0
 input [9:0] Pix_522, // sfix10_En0
 input [9:0] Pix_523, // sfix10_En0
 input [9:0] Pix_524, // sfix10_En0
 input [9:0] Pix_525, // sfix10_En0
 input [9:0] Pix_526, // sfix10_En0
 input [9:0] Pix_527, // sfix10_En0
 input [9:0] Pix_528, // sfix10_En0
 input [9:0] Pix_529, // sfix10_En0
 input [9:0] Pix_530, // sfix10_En0
 input [9:0] Pix_531, // sfix10_En0
 input [9:0] Pix_532, // sfix10_En0
 input [9:0] Pix_533, // sfix10_En0
 input [9:0] Pix_534, // sfix10_En0
 input [9:0] Pix_535, // sfix10_En0
 input [9:0] Pix_536, // sfix10_En0
 input [9:0] Pix_537, // sfix10_En0
 input [9:0] Pix_538, // sfix10_En0
 input [9:0] Pix_539, // sfix10_En0
 input [9:0] Pix_540, // sfix10_En0
 input [9:0] Pix_541, // sfix10_En0
 input [9:0] Pix_542, // sfix10_En0
 input [9:0] Pix_543, // sfix10_En0
 input [9:0] Pix_544, // sfix10_En0
 input [9:0] Pix_545, // sfix10_En0
 input [9:0] Pix_546, // sfix10_En0
 input [9:0] Pix_547, // sfix10_En0
 input [9:0] Pix_548, // sfix10_En0
 input [9:0] Pix_549, // sfix10_En0
 input [9:0] Pix_550, // sfix10_En0
 input [9:0] Pix_551, // sfix10_En0
 input [9:0] Pix_552, // sfix10_En0
 input [9:0] Pix_553, // sfix10_En0
 input [9:0] Pix_554, // sfix10_En0
 input [9:0] Pix_555, // sfix10_En0
 input [9:0] Pix_556, // sfix10_En0
 input [9:0] Pix_557, // sfix10_En0
 input [9:0] Pix_558, // sfix10_En0
 input [9:0] Pix_559, // sfix10_En0
 input [9:0] Pix_560, // sfix10_En0
 input [9:0] Pix_561, // sfix10_En0
 input [9:0] Pix_562, // sfix10_En0
 input [9:0] Pix_563, // sfix10_En0
 input [9:0] Pix_564, // sfix10_En0
 input [9:0] Pix_565, // sfix10_En0
 input [9:0] Pix_566, // sfix10_En0
 input [9:0] Pix_567, // sfix10_En0
 input [9:0] Pix_568, // sfix10_En0
 input [9:0] Pix_569, // sfix10_En0
 input [9:0] Pix_570, // sfix10_En0
 input [9:0] Pix_571, // sfix10_En0
 input [9:0] Pix_572, // sfix10_En0
 input [9:0] Pix_573, // sfix10_En0
 input [9:0] Pix_574, // sfix10_En0
 input [9:0] Pix_575, // sfix10_En0
 input [9:0] Pix_576, // sfix10_En0
 input [9:0] Pix_577, // sfix10_En0
 input [9:0] Pix_578, // sfix10_En0
 input [9:0] Pix_579, // sfix10_En0
 input [9:0] Pix_580, // sfix10_En0
 input [9:0] Pix_581, // sfix10_En0
 input [9:0] Pix_582, // sfix10_En0
 input [9:0] Pix_583, // sfix10_En0
 input [9:0] Pix_584, // sfix10_En0
 input [9:0] Pix_585, // sfix10_En0
 input [9:0] Pix_586, // sfix10_En0
 input [9:0] Pix_587, // sfix10_En0
 input [9:0] Pix_588, // sfix10_En0
 input [9:0] Pix_589, // sfix10_En0
 input [9:0] Pix_590, // sfix10_En0
 input [9:0] Pix_591, // sfix10_En0
 input [9:0] Pix_592, // sfix10_En0
 input [9:0] Pix_593, // sfix10_En0
 input [9:0] Pix_594, // sfix10_En0
 input [9:0] Pix_595, // sfix10_En0
 input [9:0] Pix_596, // sfix10_En0
 input [9:0] Pix_597, // sfix10_En0
 input [9:0] Pix_598, // sfix10_En0
 input [9:0] Pix_599, // sfix10_En0
 input [9:0] Pix_600, // sfix10_En0
 input [9:0] Pix_601, // sfix10_En0
 input [9:0] Pix_602, // sfix10_En0
 input [9:0] Pix_603, // sfix10_En0
 input [9:0] Pix_604, // sfix10_En0
 input [9:0] Pix_605, // sfix10_En0
 input [9:0] Pix_606, // sfix10_En0
 input [9:0] Pix_607, // sfix10_En0
 input [9:0] Pix_608, // sfix10_En0
 input [9:0] Pix_609, // sfix10_En0
 input [9:0] Pix_610, // sfix10_En0
 input [9:0] Pix_611, // sfix10_En0
 input [9:0] Pix_612, // sfix10_En0
 input [9:0] Pix_613, // sfix10_En0
 input [9:0] Pix_614, // sfix10_En0
 input [9:0] Pix_615, // sfix10_En0
 input [9:0] Pix_616, // sfix10_En0
 input [9:0] Pix_617, // sfix10_En0
 input [9:0] Pix_618, // sfix10_En0
 input [9:0] Pix_619, // sfix10_En0
 input [9:0] Pix_620, // sfix10_En0
 input [9:0] Pix_621, // sfix10_En0
 input [9:0] Pix_622, // sfix10_En0
 input [9:0] Pix_623, // sfix10_En0
 input [9:0] Pix_624, // sfix10_En0
 input [9:0] Pix_625, // sfix10_En0
 input [9:0] Pix_626, // sfix10_En0
 input [9:0] Pix_627, // sfix10_En0
 input [9:0] Pix_628, // sfix10_En0
 input [9:0] Pix_629, // sfix10_En0
 input [9:0] Pix_630, // sfix10_En0
 input [9:0] Pix_631, // sfix10_En0
 input [9:0] Pix_632, // sfix10_En0
 input [9:0] Pix_633, // sfix10_En0
 input [9:0] Pix_634, // sfix10_En0
 input [9:0] Pix_635, // sfix10_En0
 input [9:0] Pix_636, // sfix10_En0
 input [9:0] Pix_637, // sfix10_En0
 input [9:0] Pix_638, // sfix10_En0
 input [9:0] Pix_639, // sfix10_En0
 input [9:0] Pix_640, // sfix10_En0
 input [9:0] Pix_641, // sfix10_En0
 input [9:0] Pix_642, // sfix10_En0
 input [9:0] Pix_643, // sfix10_En0
 input [9:0] Pix_644, // sfix10_En0
 input [9:0] Pix_645, // sfix10_En0
 input [9:0] Pix_646, // sfix10_En0
 input [9:0] Pix_647, // sfix10_En0
 input [9:0] Pix_648, // sfix10_En0
 input [9:0] Pix_649, // sfix10_En0
 input [9:0] Pix_650, // sfix10_En0
 input [9:0] Pix_651, // sfix10_En0
 input [9:0] Pix_652, // sfix10_En0
 input [9:0] Pix_653, // sfix10_En0
 input [9:0] Pix_654, // sfix10_En0
 input [9:0] Pix_655, // sfix10_En0
 input [9:0] Pix_656, // sfix10_En0
 input [9:0] Pix_657, // sfix10_En0
 input [9:0] Pix_658, // sfix10_En0
 input [9:0] Pix_659, // sfix10_En0
 input [9:0] Pix_660, // sfix10_En0
 input [9:0] Pix_661, // sfix10_En0
 input [9:0] Pix_662, // sfix10_En0
 input [9:0] Pix_663, // sfix10_En0
 input [9:0] Pix_664, // sfix10_En0
 input [9:0] Pix_665, // sfix10_En0
 input [9:0] Pix_666, // sfix10_En0
 input [9:0] Pix_667, // sfix10_En0
 input [9:0] Pix_668, // sfix10_En0
 input [9:0] Pix_669, // sfix10_En0
 input [9:0] Pix_670, // sfix10_En0
 input [9:0] Pix_671, // sfix10_En0
 input [9:0] Pix_672, // sfix10_En0
 input [9:0] Pix_673, // sfix10_En0
 input [9:0] Pix_674, // sfix10_En0
 input [9:0] Pix_675, // sfix10_En0
 input [9:0] Pix_676, // sfix10_En0
 input [9:0] Pix_677, // sfix10_En0
 input [9:0] Pix_678, // sfix10_En0
 input [9:0] Pix_679, // sfix10_En0
 input [9:0] Pix_680, // sfix10_En0
 input [9:0] Pix_681, // sfix10_En0
 input [9:0] Pix_682, // sfix10_En0
 input [9:0] Pix_683, // sfix10_En0
 input [9:0] Pix_684, // sfix10_En0
 input [9:0] Pix_685, // sfix10_En0
 input [9:0] Pix_686, // sfix10_En0
 input [9:0] Pix_687, // sfix10_En0
 input [9:0] Pix_688, // sfix10_En0
 input [9:0] Pix_689, // sfix10_En0
 input [9:0] Pix_690, // sfix10_En0
 input [9:0] Pix_691, // sfix10_En0
 input [9:0] Pix_692, // sfix10_En0
 input [9:0] Pix_693, // sfix10_En0
 input [9:0] Pix_694, // sfix10_En0
 input [9:0] Pix_695, // sfix10_En0
 input [9:0] Pix_696, // sfix10_En0
 input [9:0] Pix_697, // sfix10_En0
 input [9:0] Pix_698, // sfix10_En0
 input [9:0] Pix_699, // sfix10_En0
 input [9:0] Pix_700, // sfix10_En0
 input [9:0] Pix_701, // sfix10_En0
 input [9:0] Pix_702, // sfix10_En0
 input [9:0] Pix_703, // sfix10_En0
 input [9:0] Pix_704, // sfix10_En0
 input [9:0] Pix_705, // sfix10_En0
 input [9:0] Pix_706, // sfix10_En0
 input [9:0] Pix_707, // sfix10_En0
 input [9:0] Pix_708, // sfix10_En0
 input [9:0] Pix_709, // sfix10_En0
 input [9:0] Pix_710, // sfix10_En0
 input [9:0] Pix_711, // sfix10_En0
 input [9:0] Pix_712, // sfix10_En0
 input [9:0] Pix_713, // sfix10_En0
 input [9:0] Pix_714, // sfix10_En0
 input [9:0] Pix_715, // sfix10_En0
 input [9:0] Pix_716, // sfix10_En0
 input [9:0] Pix_717, // sfix10_En0
 input [9:0] Pix_718, // sfix10_En0
 input [9:0] Pix_719, // sfix10_En0
 input [9:0] Pix_720, // sfix10_En0
 input [9:0] Pix_721, // sfix10_En0
 input [9:0] Pix_722, // sfix10_En0
 input [9:0] Pix_723, // sfix10_En0
 input [9:0] Pix_724, // sfix10_En0
 input [9:0] Pix_725, // sfix10_En0
 input [9:0] Pix_726, // sfix10_En0
 input [9:0] Pix_727, // sfix10_En0
 input [9:0] Pix_728, // sfix10_En0
 input [9:0] Pix_729, // sfix10_En0
 input [9:0] Pix_730, // sfix10_En0
 input [9:0] Pix_731, // sfix10_En0
 input [9:0] Pix_732, // sfix10_En0
 input [9:0] Pix_733, // sfix10_En0
 input [9:0] Pix_734, // sfix10_En0
 input [9:0] Pix_735, // sfix10_En0
 input [9:0] Pix_736, // sfix10_En0
 input [9:0] Pix_737, // sfix10_En0
 input [9:0] Pix_738, // sfix10_En0
 input [9:0] Pix_739, // sfix10_En0
 input [9:0] Pix_740, // sfix10_En0
 input [9:0] Pix_741, // sfix10_En0
 input [9:0] Pix_742, // sfix10_En0
 input [9:0] Pix_743, // sfix10_En0
 input [9:0] Pix_744, // sfix10_En0
 input [9:0] Pix_745, // sfix10_En0
 input [9:0] Pix_746, // sfix10_En0
 input [9:0] Pix_747, // sfix10_En0
 input [9:0] Pix_748, // sfix10_En0
 input [9:0] Pix_749, // sfix10_En0
 input [9:0] Pix_750, // sfix10_En0
 input [9:0] Pix_751, // sfix10_En0
 input [9:0] Pix_752, // sfix10_En0
 input [9:0] Pix_753, // sfix10_En0
 input [9:0] Pix_754, // sfix10_En0
 input [9:0] Pix_755, // sfix10_En0
 input [9:0] Pix_756, // sfix10_En0
 input [9:0] Pix_757, // sfix10_En0
 input [9:0] Pix_758, // sfix10_En0
 input [9:0] Pix_759, // sfix10_En0
 input [9:0] Pix_760, // sfix10_En0
 input [9:0] Pix_761, // sfix10_En0
 input [9:0] Pix_762, // sfix10_En0
 input [9:0] Pix_763, // sfix10_En0
 input [9:0] Pix_764, // sfix10_En0
 input [9:0] Pix_765, // sfix10_En0
 input [9:0] Pix_766, // sfix10_En0
 input [9:0] Pix_767, // sfix10_En0
 input [9:0] Pix_768, // sfix10_En0
 input [9:0] Pix_769, // sfix10_En0
 input [9:0] Pix_770, // sfix10_En0
 input [9:0] Pix_771, // sfix10_En0
 input [9:0] Pix_772, // sfix10_En0
 input [9:0] Pix_773, // sfix10_En0
 input [9:0] Pix_774, // sfix10_En0
 input [9:0] Pix_775, // sfix10_En0
 input [9:0] Pix_776, // sfix10_En0
 input [9:0] Pix_777, // sfix10_En0
 input [9:0] Pix_778, // sfix10_En0
 input [9:0] Pix_779, // sfix10_En0
 input [9:0] Pix_780, // sfix10_En0
 input [9:0] Pix_781, // sfix10_En0
 input [9:0] Pix_782, // sfix10_En0
 input [9:0] Pix_783, // sfix10_En0
 input [9:0] Pix_784, // sfix10_En0
 output [3:0] Image_Number, // sfix26_En18
 output reg Output_Valid
 );

// Testbench has active-low global reset
// All the blocks and modules have active-high global reset
wire globalreset;
assign globalreset = !GlobalReset;

// Set a clk to control neurons
// Input_Valid only asserts for 10 clock cycles, need another valid sign to control timing
// Multipliers and adders clk can be furthered specified to turn them off immediately when their work is done
// Not sure if this could help in power consumption
reg valid_sign;
always @(posedge clk) begin
  if(globalreset)
    valid_sign <= 0;
  else begin
    if(Input_Valid && (!Output_Valid))
	  valid_sign <= 1;
	else if(Output_Valid)
	  valid_sign <= 0;
	else
	  valid_sign <= valid_sign;
  end
end

wire neuron_clk;
assign neuron_clk = valid_sign? clk: 0;

// Timing controller
reg [9:0] N;

always @(posedge neuron_clk) begin
  if(globalreset) // Assume Input_Valid will assert til the output is ready
    N <= 0;
  else
    if(valid_sign)
      N <= N + 1;
	else
	  N <= 0;
end

// Pixel into each neurons  calvin
wire [9:0] neuron_mul_0_p, neuron_mul_1_p, neuron_mul_2_p, neuron_mul_3_p, neuron_mul_4_p, neuron_mul_5_p;
wire [9:0] neuron_mul_6_p, neuron_mul_7_p, neuron_mul_8_p, neuron_mul_9_p, neuron_mul_10_p, neuron_mul_11_p;
wire [9:0] neuron_mul_12_p, neuron_mul_13_p, neuron_mul_14_p, neuron_mul_15_p, neuron_mul_16_p, neuron_mul_17_p;
wire [9:0] neuron_mul_18_p, neuron_mul_19_p, neuron_mul_20_p, neuron_mul_21_p, neuron_mul_22_p, neuron_mul_23_p;
wire [9:0] neuron_mul_24_p, neuron_mul_25_p, neuron_mul_26_p, neuron_mul_27_p;

// Weight into each neurons
wire [18:0] neuron_0_mul_0_w, neuron_0_mul_1_w, neuron_0_mul_2_w, neuron_0_mul_3_w, neuron_0_mul_4_w, neuron_0_mul_5_w;
wire [18:0] neuron_0_mul_6_w, neuron_0_mul_7_w, neuron_0_mul_8_w, neuron_0_mul_9_w, neuron_0_mul_10_w, neuron_0_mul_11_w;
wire [18:0] neuron_0_mul_12_w, neuron_0_mul_13_w, neuron_0_mul_14_w, neuron_0_mul_15_w, neuron_0_mul_16_w, neuron_0_mul_17_w;
wire [18:0] neuron_0_mul_18_w, neuron_0_mul_19_w, neuron_0_mul_20_w, neuron_0_mul_21_w, neuron_0_mul_22_w, neuron_0_mul_23_w;
wire [18:0] neuron_0_mul_24_w, neuron_0_mul_25_w, neuron_0_mul_26_w, neuron_0_mul_27_w;

wire [18:0] neuron_1_mul_0_w, neuron_1_mul_1_w, neuron_1_mul_2_w, neuron_1_mul_3_w, neuron_1_mul_4_w, neuron_1_mul_5_w;
wire [18:0] neuron_1_mul_6_w, neuron_1_mul_7_w, neuron_1_mul_8_w, neuron_1_mul_9_w, neuron_1_mul_10_w, neuron_1_mul_11_w;
wire [18:0] neuron_1_mul_12_w, neuron_1_mul_13_w, neuron_1_mul_14_w, neuron_1_mul_15_w, neuron_1_mul_16_w, neuron_1_mul_17_w;
wire [18:0] neuron_1_mul_18_w, neuron_1_mul_19_w, neuron_1_mul_20_w, neuron_1_mul_21_w, neuron_1_mul_22_w, neuron_1_mul_23_w;
wire [18:0] neuron_1_mul_24_w, neuron_1_mul_25_w, neuron_1_mul_26_w, neuron_1_mul_27_w;

wire [18:0] neuron_2_mul_0_w, neuron_2_mul_1_w, neuron_2_mul_2_w, neuron_2_mul_3_w, neuron_2_mul_4_w, neuron_2_mul_5_w;
wire [18:0] neuron_2_mul_6_w, neuron_2_mul_7_w, neuron_2_mul_8_w, neuron_2_mul_9_w, neuron_2_mul_10_w, neuron_2_mul_11_w;
wire [18:0] neuron_2_mul_12_w, neuron_2_mul_13_w, neuron_2_mul_14_w, neuron_2_mul_15_w, neuron_2_mul_16_w, neuron_2_mul_17_w;
wire [18:0] neuron_2_mul_18_w, neuron_2_mul_19_w, neuron_2_mul_20_w, neuron_2_mul_21_w, neuron_2_mul_22_w, neuron_2_mul_23_w;
wire [18:0] neuron_2_mul_24_w, neuron_2_mul_25_w, neuron_2_mul_26_w, neuron_2_mul_27_w;

wire [18:0] neuron_3_mul_0_w, neuron_3_mul_1_w, neuron_3_mul_2_w, neuron_3_mul_3_w, neuron_3_mul_4_w, neuron_3_mul_5_w;
wire [18:0] neuron_3_mul_6_w, neuron_3_mul_7_w, neuron_3_mul_8_w, neuron_3_mul_9_w, neuron_3_mul_10_w, neuron_3_mul_11_w;
wire [18:0] neuron_3_mul_12_w, neuron_3_mul_13_w, neuron_3_mul_14_w, neuron_3_mul_15_w, neuron_3_mul_16_w, neuron_3_mul_17_w;
wire [18:0] neuron_3_mul_18_w, neuron_3_mul_19_w, neuron_3_mul_20_w, neuron_3_mul_21_w, neuron_3_mul_22_w, neuron_3_mul_23_w;
wire [18:0] neuron_3_mul_24_w, neuron_3_mul_25_w, neuron_3_mul_26_w, neuron_3_mul_27_w;

wire [18:0] neuron_4_mul_0_w, neuron_4_mul_1_w, neuron_4_mul_2_w, neuron_4_mul_3_w, neuron_4_mul_4_w, neuron_4_mul_5_w;
wire [18:0] neuron_4_mul_6_w, neuron_4_mul_7_w, neuron_4_mul_8_w, neuron_4_mul_9_w, neuron_4_mul_10_w, neuron_4_mul_11_w;
wire [18:0] neuron_4_mul_12_w, neuron_4_mul_13_w, neuron_4_mul_14_w, neuron_4_mul_15_w, neuron_4_mul_16_w, neuron_4_mul_17_w;
wire [18:0] neuron_4_mul_18_w, neuron_4_mul_19_w, neuron_4_mul_20_w, neuron_4_mul_21_w, neuron_4_mul_22_w, neuron_4_mul_23_w;
wire [18:0] neuron_4_mul_24_w, neuron_4_mul_25_w, neuron_4_mul_26_w, neuron_4_mul_27_w;

wire [18:0] neuron_5_mul_0_w, neuron_5_mul_1_w, neuron_5_mul_2_w, neuron_5_mul_3_w, neuron_5_mul_4_w, neuron_5_mul_5_w;
wire [18:0] neuron_5_mul_6_w, neuron_5_mul_7_w, neuron_5_mul_8_w, neuron_5_mul_9_w, neuron_5_mul_10_w, neuron_5_mul_11_w;
wire [18:0] neuron_5_mul_12_w, neuron_5_mul_13_w, neuron_5_mul_14_w, neuron_5_mul_15_w, neuron_5_mul_16_w, neuron_5_mul_17_w;
wire [18:0] neuron_5_mul_18_w, neuron_5_mul_19_w, neuron_5_mul_20_w, neuron_5_mul_21_w, neuron_5_mul_22_w, neuron_5_mul_23_w;
wire [18:0] neuron_5_mul_24_w, neuron_5_mul_25_w, neuron_5_mul_26_w, neuron_5_mul_27_w;

wire [18:0] neuron_6_mul_0_w, neuron_6_mul_1_w, neuron_6_mul_2_w, neuron_6_mul_3_w, neuron_6_mul_4_w, neuron_6_mul_5_w;
wire [18:0] neuron_6_mul_6_w, neuron_6_mul_7_w, neuron_6_mul_8_w, neuron_6_mul_9_w, neuron_6_mul_10_w, neuron_6_mul_11_w;
wire [18:0] neuron_6_mul_12_w, neuron_6_mul_13_w, neuron_6_mul_14_w, neuron_6_mul_15_w, neuron_6_mul_16_w, neuron_6_mul_17_w;
wire [18:0] neuron_6_mul_18_w, neuron_6_mul_19_w, neuron_6_mul_20_w, neuron_6_mul_21_w, neuron_6_mul_22_w, neuron_6_mul_23_w;
wire [18:0] neuron_6_mul_24_w, neuron_6_mul_25_w, neuron_6_mul_26_w, neuron_6_mul_27_w;

wire [18:0] neuron_7_mul_0_w, neuron_7_mul_1_w, neuron_7_mul_2_w, neuron_7_mul_3_w, neuron_7_mul_4_w, neuron_7_mul_5_w;
wire [18:0] neuron_7_mul_6_w, neuron_7_mul_7_w, neuron_7_mul_8_w, neuron_7_mul_9_w, neuron_7_mul_10_w, neuron_7_mul_11_w;
wire [18:0] neuron_7_mul_12_w, neuron_7_mul_13_w, neuron_7_mul_14_w, neuron_7_mul_15_w, neuron_7_mul_16_w, neuron_7_mul_17_w;
wire [18:0] neuron_7_mul_18_w, neuron_7_mul_19_w, neuron_7_mul_20_w, neuron_7_mul_21_w, neuron_7_mul_22_w, neuron_7_mul_23_w;
wire [18:0] neuron_7_mul_24_w, neuron_7_mul_25_w, neuron_7_mul_26_w, neuron_7_mul_27_w;

wire [18:0] neuron_8_mul_0_w, neuron_8_mul_1_w, neuron_8_mul_2_w, neuron_8_mul_3_w, neuron_8_mul_4_w, neuron_8_mul_5_w;
wire [18:0] neuron_8_mul_6_w, neuron_8_mul_7_w, neuron_8_mul_8_w, neuron_8_mul_9_w, neuron_8_mul_10_w, neuron_8_mul_11_w;
wire [18:0] neuron_8_mul_12_w, neuron_8_mul_13_w, neuron_8_mul_14_w, neuron_8_mul_15_w, neuron_8_mul_16_w, neuron_8_mul_17_w;
wire [18:0] neuron_8_mul_18_w, neuron_8_mul_19_w, neuron_8_mul_20_w, neuron_8_mul_21_w, neuron_8_mul_22_w, neuron_8_mul_23_w;
wire [18:0] neuron_8_mul_24_w, neuron_8_mul_25_w, neuron_8_mul_26_w, neuron_8_mul_27_w;

wire [18:0] neuron_9_mul_0_w, neuron_9_mul_1_w, neuron_9_mul_2_w, neuron_9_mul_3_w, neuron_9_mul_4_w, neuron_9_mul_5_w;
wire [18:0] neuron_9_mul_6_w, neuron_9_mul_7_w, neuron_9_mul_8_w, neuron_9_mul_9_w, neuron_9_mul_10_w, neuron_9_mul_11_w;
wire [18:0] neuron_9_mul_12_w, neuron_9_mul_13_w, neuron_9_mul_14_w, neuron_9_mul_15_w, neuron_9_mul_16_w, neuron_9_mul_17_w;
wire [18:0] neuron_9_mul_18_w, neuron_9_mul_19_w, neuron_9_mul_20_w, neuron_9_mul_21_w, neuron_9_mul_22_w, neuron_9_mul_23_w;
wire [18:0] neuron_9_mul_24_w, neuron_9_mul_25_w, neuron_9_mul_26_w, neuron_9_mul_27_w;

// Output of each multiplier 28*10
wire [25:0] neuron_0_mul_0_out, neuron_0_mul_1_out, neuron_0_mul_2_out, neuron_0_mul_3_out, neuron_0_mul_4_out;
wire [25:0] neuron_0_mul_5_out, neuron_0_mul_6_out, neuron_0_mul_7_out, neuron_0_mul_8_out, neuron_0_mul_9_out;
wire [25:0] neuron_0_mul_10_out, neuron_0_mul_11_out, neuron_0_mul_12_out, neuron_0_mul_13_out, neuron_0_mul_14_out;
wire [25:0] neuron_0_mul_15_out, neuron_0_mul_16_out, neuron_0_mul_17_out, neuron_0_mul_18_out, neuron_0_mul_19_out;
wire [25:0] neuron_0_mul_20_out, neuron_0_mul_21_out, neuron_0_mul_22_out, neuron_0_mul_23_out, neuron_0_mul_24_out;
wire [25:0] neuron_0_mul_25_out, neuron_0_mul_26_out, neuron_0_mul_27_out;

wire [25:0] neuron_1_mul_0_out, neuron_1_mul_1_out, neuron_1_mul_2_out, neuron_1_mul_3_out, neuron_1_mul_4_out;
wire [25:0] neuron_1_mul_5_out, neuron_1_mul_6_out, neuron_1_mul_7_out, neuron_1_mul_8_out, neuron_1_mul_9_out;
wire [25:0] neuron_1_mul_10_out, neuron_1_mul_11_out, neuron_1_mul_12_out, neuron_1_mul_13_out, neuron_1_mul_14_out;
wire [25:0] neuron_1_mul_15_out, neuron_1_mul_16_out, neuron_1_mul_17_out, neuron_1_mul_18_out, neuron_1_mul_19_out;
wire [25:0] neuron_1_mul_20_out, neuron_1_mul_21_out, neuron_1_mul_22_out, neuron_1_mul_23_out, neuron_1_mul_24_out;
wire [25:0] neuron_1_mul_25_out, neuron_1_mul_26_out, neuron_1_mul_27_out;

wire [25:0] neuron_2_mul_0_out, neuron_2_mul_1_out, neuron_2_mul_2_out, neuron_2_mul_3_out, neuron_2_mul_4_out;
wire [25:0] neuron_2_mul_5_out, neuron_2_mul_6_out, neuron_2_mul_7_out, neuron_2_mul_8_out, neuron_2_mul_9_out;
wire [25:0] neuron_2_mul_10_out, neuron_2_mul_11_out, neuron_2_mul_12_out, neuron_2_mul_13_out, neuron_2_mul_14_out;
wire [25:0] neuron_2_mul_15_out, neuron_2_mul_16_out, neuron_2_mul_17_out, neuron_2_mul_18_out, neuron_2_mul_19_out;
wire [25:0] neuron_2_mul_20_out, neuron_2_mul_21_out, neuron_2_mul_22_out, neuron_2_mul_23_out, neuron_2_mul_24_out;
wire [25:0] neuron_2_mul_25_out, neuron_2_mul_26_out, neuron_2_mul_27_out;

wire [25:0] neuron_3_mul_0_out, neuron_3_mul_1_out, neuron_3_mul_2_out, neuron_3_mul_3_out, neuron_3_mul_4_out;
wire [25:0] neuron_3_mul_5_out, neuron_3_mul_6_out, neuron_3_mul_7_out, neuron_3_mul_8_out, neuron_3_mul_9_out;
wire [25:0] neuron_3_mul_10_out, neuron_3_mul_11_out, neuron_3_mul_12_out, neuron_3_mul_13_out, neuron_3_mul_14_out;
wire [25:0] neuron_3_mul_15_out, neuron_3_mul_16_out, neuron_3_mul_17_out, neuron_3_mul_18_out, neuron_3_mul_19_out;
wire [25:0] neuron_3_mul_20_out, neuron_3_mul_21_out, neuron_3_mul_22_out, neuron_3_mul_23_out, neuron_3_mul_24_out;
wire [25:0] neuron_3_mul_25_out, neuron_3_mul_26_out, neuron_3_mul_27_out;

wire [25:0] neuron_4_mul_0_out, neuron_4_mul_1_out, neuron_4_mul_2_out, neuron_4_mul_3_out, neuron_4_mul_4_out;
wire [25:0] neuron_4_mul_5_out, neuron_4_mul_6_out, neuron_4_mul_7_out, neuron_4_mul_8_out, neuron_4_mul_9_out;
wire [25:0] neuron_4_mul_10_out, neuron_4_mul_11_out, neuron_4_mul_12_out, neuron_4_mul_13_out, neuron_4_mul_14_out;
wire [25:0] neuron_4_mul_15_out, neuron_4_mul_16_out, neuron_4_mul_17_out, neuron_4_mul_18_out, neuron_4_mul_19_out;
wire [25:0] neuron_4_mul_20_out, neuron_4_mul_21_out, neuron_4_mul_22_out, neuron_4_mul_23_out, neuron_4_mul_24_out;
wire [25:0] neuron_4_mul_25_out, neuron_4_mul_26_out, neuron_4_mul_27_out;

wire [25:0] neuron_5_mul_0_out, neuron_5_mul_1_out, neuron_5_mul_2_out, neuron_5_mul_3_out, neuron_5_mul_4_out;
wire [25:0] neuron_5_mul_5_out, neuron_5_mul_6_out, neuron_5_mul_7_out, neuron_5_mul_8_out, neuron_5_mul_9_out;
wire [25:0] neuron_5_mul_10_out, neuron_5_mul_11_out, neuron_5_mul_12_out, neuron_5_mul_13_out, neuron_5_mul_14_out;
wire [25:0] neuron_5_mul_15_out, neuron_5_mul_16_out, neuron_5_mul_17_out, neuron_5_mul_18_out, neuron_5_mul_19_out;
wire [25:0] neuron_5_mul_20_out, neuron_5_mul_21_out, neuron_5_mul_22_out, neuron_5_mul_23_out, neuron_5_mul_24_out;
wire [25:0] neuron_5_mul_25_out, neuron_5_mul_26_out, neuron_5_mul_27_out;

wire [25:0] neuron_6_mul_0_out, neuron_6_mul_1_out, neuron_6_mul_2_out, neuron_6_mul_3_out, neuron_6_mul_4_out;
wire [25:0] neuron_6_mul_5_out, neuron_6_mul_6_out, neuron_6_mul_7_out, neuron_6_mul_8_out, neuron_6_mul_9_out;
wire [25:0] neuron_6_mul_10_out, neuron_6_mul_11_out, neuron_6_mul_12_out, neuron_6_mul_13_out, neuron_6_mul_14_out;
wire [25:0] neuron_6_mul_15_out, neuron_6_mul_16_out, neuron_6_mul_17_out, neuron_6_mul_18_out, neuron_6_mul_19_out;
wire [25:0] neuron_6_mul_20_out, neuron_6_mul_21_out, neuron_6_mul_22_out, neuron_6_mul_23_out, neuron_6_mul_24_out;
wire [25:0] neuron_6_mul_25_out, neuron_6_mul_26_out, neuron_6_mul_27_out;

wire [25:0] neuron_7_mul_0_out, neuron_7_mul_1_out, neuron_7_mul_2_out, neuron_7_mul_3_out, neuron_7_mul_4_out;
wire [25:0] neuron_7_mul_5_out, neuron_7_mul_6_out, neuron_7_mul_7_out, neuron_7_mul_8_out, neuron_7_mul_9_out;
wire [25:0] neuron_7_mul_10_out, neuron_7_mul_11_out, neuron_7_mul_12_out, neuron_7_mul_13_out, neuron_7_mul_14_out;
wire [25:0] neuron_7_mul_15_out, neuron_7_mul_16_out, neuron_7_mul_17_out, neuron_7_mul_18_out, neuron_7_mul_19_out;
wire [25:0] neuron_7_mul_20_out, neuron_7_mul_21_out, neuron_7_mul_22_out, neuron_7_mul_23_out, neuron_7_mul_24_out;
wire [25:0] neuron_7_mul_25_out, neuron_7_mul_26_out, neuron_7_mul_27_out;

wire [25:0] neuron_8_mul_0_out, neuron_8_mul_1_out, neuron_8_mul_2_out, neuron_8_mul_3_out, neuron_8_mul_4_out;
wire [25:0] neuron_8_mul_5_out, neuron_8_mul_6_out, neuron_8_mul_7_out, neuron_8_mul_8_out, neuron_8_mul_9_out;
wire [25:0] neuron_8_mul_10_out, neuron_8_mul_11_out, neuron_8_mul_12_out, neuron_8_mul_13_out, neuron_8_mul_14_out;
wire [25:0] neuron_8_mul_15_out, neuron_8_mul_16_out, neuron_8_mul_17_out, neuron_8_mul_18_out, neuron_8_mul_19_out;
wire [25:0] neuron_8_mul_20_out, neuron_8_mul_21_out, neuron_8_mul_22_out, neuron_8_mul_23_out, neuron_8_mul_24_out;
wire [25:0] neuron_8_mul_25_out, neuron_8_mul_26_out, neuron_8_mul_27_out;

wire [25:0] neuron_9_mul_0_out, neuron_9_mul_1_out, neuron_9_mul_2_out, neuron_9_mul_3_out, neuron_9_mul_4_out;
wire [25:0] neuron_9_mul_5_out, neuron_9_mul_6_out, neuron_9_mul_7_out, neuron_9_mul_8_out, neuron_9_mul_9_out;
wire [25:0] neuron_9_mul_10_out, neuron_9_mul_11_out, neuron_9_mul_12_out, neuron_9_mul_13_out, neuron_9_mul_14_out;
wire [25:0] neuron_9_mul_15_out, neuron_9_mul_16_out, neuron_9_mul_17_out, neuron_9_mul_18_out, neuron_9_mul_19_out;
wire [25:0] neuron_9_mul_20_out, neuron_9_mul_21_out, neuron_9_mul_22_out, neuron_9_mul_23_out, neuron_9_mul_24_out;
wire [25:0] neuron_9_mul_25_out, neuron_9_mul_26_out, neuron_9_mul_27_out;



// Input number of each adder 28*10
wire [25:0] neuron_0_add_0_p1, neuron_0_add_0_p2, neuron_0_add_1_p1, neuron_0_add_1_p2, neuron_0_add_2_p1, neuron_0_add_2_p2, neuron_0_add_3_p1, neuron_0_add_3_p2;
wire [25:0] neuron_0_add_4_p1, neuron_0_add_4_p2, neuron_0_add_5_p1, neuron_0_add_5_p2, neuron_0_add_6_p1, neuron_0_add_6_p2, neuron_0_add_7_p1, neuron_0_add_7_p2;
wire [25:0] neuron_0_add_8_p1, neuron_0_add_8_p2, neuron_0_add_9_p1, neuron_0_add_9_p2, neuron_0_add_10_p1, neuron_0_add_10_p2, neuron_0_add_11_p1, neuron_0_add_11_p2;
wire [25:0] neuron_0_add_12_p1, neuron_0_add_12_p2, neuron_0_add_13_p1, neuron_0_add_13_p2, neuron_0_add_14_p1, neuron_0_add_14_p2, neuron_0_add_15_p1, neuron_0_add_15_p2;
wire [25:0] neuron_0_add_16_p1, neuron_0_add_16_p2, neuron_0_add_17_p1, neuron_0_add_17_p2, neuron_0_add_18_p1, neuron_0_add_18_p2, neuron_0_add_19_p1, neuron_0_add_19_p2;
wire [25:0] neuron_0_add_20_p1, neuron_0_add_20_p2, neuron_0_add_21_p1, neuron_0_add_21_p2, neuron_0_add_22_p1, neuron_0_add_22_p2, neuron_0_add_23_p1, neuron_0_add_23_p2;
wire [25:0] neuron_0_add_24_p1, neuron_0_add_24_p2, neuron_0_add_25_p1, neuron_0_add_25_p2, neuron_0_add_26_p1, neuron_0_add_26_p2, neuron_0_add_27_p1, neuron_0_add_27_p2;

wire [25:0] neuron_1_add_0_p1, neuron_1_add_0_p2, neuron_1_add_1_p1, neuron_1_add_1_p2, neuron_1_add_2_p1, neuron_1_add_2_p2, neuron_1_add_3_p1, neuron_1_add_3_p2;
wire [25:0] neuron_1_add_4_p1, neuron_1_add_4_p2, neuron_1_add_5_p1, neuron_1_add_5_p2, neuron_1_add_6_p1, neuron_1_add_6_p2, neuron_1_add_7_p1, neuron_1_add_7_p2;
wire [25:0] neuron_1_add_8_p1, neuron_1_add_8_p2, neuron_1_add_9_p1, neuron_1_add_9_p2, neuron_1_add_10_p1, neuron_1_add_10_p2, neuron_1_add_11_p1, neuron_1_add_11_p2;
wire [25:0] neuron_1_add_12_p1, neuron_1_add_12_p2, neuron_1_add_13_p1, neuron_1_add_13_p2, neuron_1_add_14_p1, neuron_1_add_14_p2, neuron_1_add_15_p1, neuron_1_add_15_p2;
wire [25:0] neuron_1_add_16_p1, neuron_1_add_16_p2, neuron_1_add_17_p1, neuron_1_add_17_p2, neuron_1_add_18_p1, neuron_1_add_18_p2, neuron_1_add_19_p1, neuron_1_add_19_p2;
wire [25:0] neuron_1_add_20_p1, neuron_1_add_20_p2, neuron_1_add_21_p1, neuron_1_add_21_p2, neuron_1_add_22_p1, neuron_1_add_22_p2, neuron_1_add_23_p1, neuron_1_add_23_p2;
wire [25:0] neuron_1_add_24_p1, neuron_1_add_24_p2, neuron_1_add_25_p1, neuron_1_add_25_p2, neuron_1_add_26_p1, neuron_1_add_26_p2, neuron_1_add_27_p1, neuron_1_add_27_p2;

wire [25:0] neuron_2_add_0_p1, neuron_2_add_0_p2, neuron_2_add_1_p1, neuron_2_add_1_p2, neuron_2_add_2_p1, neuron_2_add_2_p2, neuron_2_add_3_p1, neuron_2_add_3_p2;
wire [25:0] neuron_2_add_4_p1, neuron_2_add_4_p2, neuron_2_add_5_p1, neuron_2_add_5_p2, neuron_2_add_6_p1, neuron_2_add_6_p2, neuron_2_add_7_p1, neuron_2_add_7_p2;
wire [25:0] neuron_2_add_8_p1, neuron_2_add_8_p2, neuron_2_add_9_p1, neuron_2_add_9_p2, neuron_2_add_10_p1, neuron_2_add_10_p2, neuron_2_add_11_p1, neuron_2_add_11_p2;
wire [25:0] neuron_2_add_12_p1, neuron_2_add_12_p2, neuron_2_add_13_p1, neuron_2_add_13_p2, neuron_2_add_14_p1, neuron_2_add_14_p2, neuron_2_add_15_p1, neuron_2_add_15_p2;
wire [25:0] neuron_2_add_16_p1, neuron_2_add_16_p2, neuron_2_add_17_p1, neuron_2_add_17_p2, neuron_2_add_18_p1, neuron_2_add_18_p2, neuron_2_add_19_p1, neuron_2_add_19_p2;
wire [25:0] neuron_2_add_20_p1, neuron_2_add_20_p2, neuron_2_add_21_p1, neuron_2_add_21_p2, neuron_2_add_22_p1, neuron_2_add_22_p2, neuron_2_add_23_p1, neuron_2_add_23_p2;
wire [25:0] neuron_2_add_24_p1, neuron_2_add_24_p2, neuron_2_add_25_p1, neuron_2_add_25_p2, neuron_2_add_26_p1, neuron_2_add_26_p2, neuron_2_add_27_p1, neuron_2_add_27_p2;

wire [25:0] neuron_3_add_0_p1, neuron_3_add_0_p2, neuron_3_add_1_p1, neuron_3_add_1_p2, neuron_3_add_2_p1, neuron_3_add_2_p2, neuron_3_add_3_p1, neuron_3_add_3_p2;
wire [25:0] neuron_3_add_4_p1, neuron_3_add_4_p2, neuron_3_add_5_p1, neuron_3_add_5_p2, neuron_3_add_6_p1, neuron_3_add_6_p2, neuron_3_add_7_p1, neuron_3_add_7_p2;
wire [25:0] neuron_3_add_8_p1, neuron_3_add_8_p2, neuron_3_add_9_p1, neuron_3_add_9_p2, neuron_3_add_10_p1, neuron_3_add_10_p2, neuron_3_add_11_p1, neuron_3_add_11_p2;
wire [25:0] neuron_3_add_12_p1, neuron_3_add_12_p2, neuron_3_add_13_p1, neuron_3_add_13_p2, neuron_3_add_14_p1, neuron_3_add_14_p2, neuron_3_add_15_p1, neuron_3_add_15_p2;
wire [25:0] neuron_3_add_16_p1, neuron_3_add_16_p2, neuron_3_add_17_p1, neuron_3_add_17_p2, neuron_3_add_18_p1, neuron_3_add_18_p2, neuron_3_add_19_p1, neuron_3_add_19_p2;
wire [25:0] neuron_3_add_20_p1, neuron_3_add_20_p2, neuron_3_add_21_p1, neuron_3_add_21_p2, neuron_3_add_22_p1, neuron_3_add_22_p2, neuron_3_add_23_p1, neuron_3_add_23_p2;
wire [25:0] neuron_3_add_24_p1, neuron_3_add_24_p2, neuron_3_add_25_p1, neuron_3_add_25_p2, neuron_3_add_26_p1, neuron_3_add_26_p2, neuron_3_add_27_p1, neuron_3_add_27_p2;

wire [25:0] neuron_4_add_0_p1, neuron_4_add_0_p2, neuron_4_add_1_p1, neuron_4_add_1_p2, neuron_4_add_2_p1, neuron_4_add_2_p2, neuron_4_add_3_p1, neuron_4_add_3_p2;
wire [25:0] neuron_4_add_4_p1, neuron_4_add_4_p2, neuron_4_add_5_p1, neuron_4_add_5_p2, neuron_4_add_6_p1, neuron_4_add_6_p2, neuron_4_add_7_p1, neuron_4_add_7_p2;
wire [25:0] neuron_4_add_8_p1, neuron_4_add_8_p2, neuron_4_add_9_p1, neuron_4_add_9_p2, neuron_4_add_10_p1, neuron_4_add_10_p2, neuron_4_add_11_p1, neuron_4_add_11_p2;
wire [25:0] neuron_4_add_12_p1, neuron_4_add_12_p2, neuron_4_add_13_p1, neuron_4_add_13_p2, neuron_4_add_14_p1, neuron_4_add_14_p2, neuron_4_add_15_p1, neuron_4_add_15_p2;
wire [25:0] neuron_4_add_16_p1, neuron_4_add_16_p2, neuron_4_add_17_p1, neuron_4_add_17_p2, neuron_4_add_18_p1, neuron_4_add_18_p2, neuron_4_add_19_p1, neuron_4_add_19_p2;
wire [25:0] neuron_4_add_20_p1, neuron_4_add_20_p2, neuron_4_add_21_p1, neuron_4_add_21_p2, neuron_4_add_22_p1, neuron_4_add_22_p2, neuron_4_add_23_p1, neuron_4_add_23_p2;
wire [25:0] neuron_4_add_24_p1, neuron_4_add_24_p2, neuron_4_add_25_p1, neuron_4_add_25_p2, neuron_4_add_26_p1, neuron_4_add_26_p2, neuron_4_add_27_p1, neuron_4_add_27_p2;

wire [25:0] neuron_5_add_0_p1, neuron_5_add_0_p2, neuron_5_add_1_p1, neuron_5_add_1_p2, neuron_5_add_2_p1, neuron_5_add_2_p2, neuron_5_add_3_p1, neuron_5_add_3_p2;
wire [25:0] neuron_5_add_4_p1, neuron_5_add_4_p2, neuron_5_add_5_p1, neuron_5_add_5_p2, neuron_5_add_6_p1, neuron_5_add_6_p2, neuron_5_add_7_p1, neuron_5_add_7_p2;
wire [25:0] neuron_5_add_8_p1, neuron_5_add_8_p2, neuron_5_add_9_p1, neuron_5_add_9_p2, neuron_5_add_10_p1, neuron_5_add_10_p2, neuron_5_add_11_p1, neuron_5_add_11_p2;
wire [25:0] neuron_5_add_12_p1, neuron_5_add_12_p2, neuron_5_add_13_p1, neuron_5_add_13_p2, neuron_5_add_14_p1, neuron_5_add_14_p2, neuron_5_add_15_p1, neuron_5_add_15_p2;
wire [25:0] neuron_5_add_16_p1, neuron_5_add_16_p2, neuron_5_add_17_p1, neuron_5_add_17_p2, neuron_5_add_18_p1, neuron_5_add_18_p2, neuron_5_add_19_p1, neuron_5_add_19_p2;
wire [25:0] neuron_5_add_20_p1, neuron_5_add_20_p2, neuron_5_add_21_p1, neuron_5_add_21_p2, neuron_5_add_22_p1, neuron_5_add_22_p2, neuron_5_add_23_p1, neuron_5_add_23_p2;
wire [25:0] neuron_5_add_24_p1, neuron_5_add_24_p2, neuron_5_add_25_p1, neuron_5_add_25_p2, neuron_5_add_26_p1, neuron_5_add_26_p2, neuron_5_add_27_p1, neuron_5_add_27_p2;

wire [25:0] neuron_6_add_0_p1, neuron_6_add_0_p2, neuron_6_add_1_p1, neuron_6_add_1_p2, neuron_6_add_2_p1, neuron_6_add_2_p2, neuron_6_add_3_p1, neuron_6_add_3_p2;
wire [25:0] neuron_6_add_4_p1, neuron_6_add_4_p2, neuron_6_add_5_p1, neuron_6_add_5_p2, neuron_6_add_6_p1, neuron_6_add_6_p2, neuron_6_add_7_p1, neuron_6_add_7_p2;
wire [25:0] neuron_6_add_8_p1, neuron_6_add_8_p2, neuron_6_add_9_p1, neuron_6_add_9_p2, neuron_6_add_10_p1, neuron_6_add_10_p2, neuron_6_add_11_p1, neuron_6_add_11_p2;
wire [25:0] neuron_6_add_12_p1, neuron_6_add_12_p2, neuron_6_add_13_p1, neuron_6_add_13_p2, neuron_6_add_14_p1, neuron_6_add_14_p2, neuron_6_add_15_p1, neuron_6_add_15_p2;
wire [25:0] neuron_6_add_16_p1, neuron_6_add_16_p2, neuron_6_add_17_p1, neuron_6_add_17_p2, neuron_6_add_18_p1, neuron_6_add_18_p2, neuron_6_add_19_p1, neuron_6_add_19_p2;
wire [25:0] neuron_6_add_20_p1, neuron_6_add_20_p2, neuron_6_add_21_p1, neuron_6_add_21_p2, neuron_6_add_22_p1, neuron_6_add_22_p2, neuron_6_add_23_p1, neuron_6_add_23_p2;
wire [25:0] neuron_6_add_24_p1, neuron_6_add_24_p2, neuron_6_add_25_p1, neuron_6_add_25_p2, neuron_6_add_26_p1, neuron_6_add_26_p2, neuron_6_add_27_p1, neuron_6_add_27_p2;

wire [25:0] neuron_7_add_0_p1, neuron_7_add_0_p2, neuron_7_add_1_p1, neuron_7_add_1_p2, neuron_7_add_2_p1, neuron_7_add_2_p2, neuron_7_add_3_p1, neuron_7_add_3_p2;
wire [25:0] neuron_7_add_4_p1, neuron_7_add_4_p2, neuron_7_add_5_p1, neuron_7_add_5_p2, neuron_7_add_6_p1, neuron_7_add_6_p2, neuron_7_add_7_p1, neuron_7_add_7_p2;
wire [25:0] neuron_7_add_8_p1, neuron_7_add_8_p2, neuron_7_add_9_p1, neuron_7_add_9_p2, neuron_7_add_10_p1, neuron_7_add_10_p2, neuron_7_add_11_p1, neuron_7_add_11_p2;
wire [25:0] neuron_7_add_12_p1, neuron_7_add_12_p2, neuron_7_add_13_p1, neuron_7_add_13_p2, neuron_7_add_14_p1, neuron_7_add_14_p2, neuron_7_add_15_p1, neuron_7_add_15_p2;
wire [25:0] neuron_7_add_16_p1, neuron_7_add_16_p2, neuron_7_add_17_p1, neuron_7_add_17_p2, neuron_7_add_18_p1, neuron_7_add_18_p2, neuron_7_add_19_p1, neuron_7_add_19_p2;
wire [25:0] neuron_7_add_20_p1, neuron_7_add_20_p2, neuron_7_add_21_p1, neuron_7_add_21_p2, neuron_7_add_22_p1, neuron_7_add_22_p2, neuron_7_add_23_p1, neuron_7_add_23_p2;
wire [25:0] neuron_7_add_24_p1, neuron_7_add_24_p2, neuron_7_add_25_p1, neuron_7_add_25_p2, neuron_7_add_26_p1, neuron_7_add_26_p2, neuron_7_add_27_p1, neuron_7_add_27_p2;

wire [25:0] neuron_8_add_0_p1, neuron_8_add_0_p2, neuron_8_add_1_p1, neuron_8_add_1_p2, neuron_8_add_2_p1, neuron_8_add_2_p2, neuron_8_add_3_p1, neuron_8_add_3_p2;
wire [25:0] neuron_8_add_4_p1, neuron_8_add_4_p2, neuron_8_add_5_p1, neuron_8_add_5_p2, neuron_8_add_6_p1, neuron_8_add_6_p2, neuron_8_add_7_p1, neuron_8_add_7_p2;
wire [25:0] neuron_8_add_8_p1, neuron_8_add_8_p2, neuron_8_add_9_p1, neuron_8_add_9_p2, neuron_8_add_10_p1, neuron_8_add_10_p2, neuron_8_add_11_p1, neuron_8_add_11_p2;
wire [25:0] neuron_8_add_12_p1, neuron_8_add_12_p2, neuron_8_add_13_p1, neuron_8_add_13_p2, neuron_8_add_14_p1, neuron_8_add_14_p2, neuron_8_add_15_p1, neuron_8_add_15_p2;
wire [25:0] neuron_8_add_16_p1, neuron_8_add_16_p2, neuron_8_add_17_p1, neuron_8_add_17_p2, neuron_8_add_18_p1, neuron_8_add_18_p2, neuron_8_add_19_p1, neuron_8_add_19_p2;
wire [25:0] neuron_8_add_20_p1, neuron_8_add_20_p2, neuron_8_add_21_p1, neuron_8_add_21_p2, neuron_8_add_22_p1, neuron_8_add_22_p2, neuron_8_add_23_p1, neuron_8_add_23_p2;
wire [25:0] neuron_8_add_24_p1, neuron_8_add_24_p2, neuron_8_add_25_p1, neuron_8_add_25_p2, neuron_8_add_26_p1, neuron_8_add_26_p2, neuron_8_add_27_p1, neuron_8_add_27_p2;

wire [25:0] neuron_9_add_0_p1, neuron_9_add_0_p2, neuron_9_add_1_p1, neuron_9_add_1_p2, neuron_9_add_2_p1, neuron_9_add_2_p2, neuron_9_add_3_p1, neuron_9_add_3_p2;
wire [25:0] neuron_9_add_4_p1, neuron_9_add_4_p2, neuron_9_add_5_p1, neuron_9_add_5_p2, neuron_9_add_6_p1, neuron_9_add_6_p2, neuron_9_add_7_p1, neuron_9_add_7_p2;
wire [25:0] neuron_9_add_8_p1, neuron_9_add_8_p2, neuron_9_add_9_p1, neuron_9_add_9_p2, neuron_9_add_10_p1, neuron_9_add_10_p2, neuron_9_add_11_p1, neuron_9_add_11_p2;
wire [25:0] neuron_9_add_12_p1, neuron_9_add_12_p2, neuron_9_add_13_p1, neuron_9_add_13_p2, neuron_9_add_14_p1, neuron_9_add_14_p2, neuron_9_add_15_p1, neuron_9_add_15_p2;
wire [25:0] neuron_9_add_16_p1, neuron_9_add_16_p2, neuron_9_add_17_p1, neuron_9_add_17_p2, neuron_9_add_18_p1, neuron_9_add_18_p2, neuron_9_add_19_p1, neuron_9_add_19_p2;
wire [25:0] neuron_9_add_20_p1, neuron_9_add_20_p2, neuron_9_add_21_p1, neuron_9_add_21_p2, neuron_9_add_22_p1, neuron_9_add_22_p2, neuron_9_add_23_p1, neuron_9_add_23_p2;
wire [25:0] neuron_9_add_24_p1, neuron_9_add_24_p2, neuron_9_add_25_p1, neuron_9_add_25_p2, neuron_9_add_26_p1, neuron_9_add_26_p2, neuron_9_add_27_p1, neuron_9_add_27_p2;

// Output of each adder
wire [25:0] neuron_0_add_0_out, neuron_0_add_1_out, neuron_0_add_2_out, neuron_0_add_3_out, neuron_0_add_4_out, neuron_0_add_5_out;
wire [25:0] neuron_0_add_6_out, neuron_0_add_7_out, neuron_0_add_8_out, neuron_0_add_9_out, neuron_0_add_10_out, neuron_0_add_11_out;
wire [25:0] neuron_0_add_12_out, neuron_0_add_13_out, neuron_0_add_14_out, neuron_0_add_15_out, neuron_0_add_16_out, neuron_0_add_17_out;
wire [25:0] neuron_0_add_18_out, neuron_0_add_19_out, neuron_0_add_20_out, neuron_0_add_21_out, neuron_0_add_22_out, neuron_0_add_23_out;
wire [25:0] neuron_0_add_24_out, neuron_0_add_25_out, neuron_0_add_26_out, neuron_0_add_27_out;

wire [25:0] neuron_1_add_0_out, neuron_1_add_1_out, neuron_1_add_2_out, neuron_1_add_3_out, neuron_1_add_4_out, neuron_1_add_5_out;
wire [25:0] neuron_1_add_6_out, neuron_1_add_7_out, neuron_1_add_8_out, neuron_1_add_9_out, neuron_1_add_10_out, neuron_1_add_11_out;
wire [25:0] neuron_1_add_12_out, neuron_1_add_13_out, neuron_1_add_14_out, neuron_1_add_15_out, neuron_1_add_16_out, neuron_1_add_17_out;
wire [25:0] neuron_1_add_18_out, neuron_1_add_19_out, neuron_1_add_20_out, neuron_1_add_21_out, neuron_1_add_22_out, neuron_1_add_23_out;
wire [25:0] neuron_1_add_24_out, neuron_1_add_25_out, neuron_1_add_26_out, neuron_1_add_27_out;

wire [25:0] neuron_2_add_0_out, neuron_2_add_1_out, neuron_2_add_2_out, neuron_2_add_3_out, neuron_2_add_4_out, neuron_2_add_5_out;
wire [25:0] neuron_2_add_6_out, neuron_2_add_7_out, neuron_2_add_8_out, neuron_2_add_9_out, neuron_2_add_10_out, neuron_2_add_11_out;
wire [25:0] neuron_2_add_12_out, neuron_2_add_13_out, neuron_2_add_14_out, neuron_2_add_15_out, neuron_2_add_16_out, neuron_2_add_17_out;
wire [25:0] neuron_2_add_18_out, neuron_2_add_19_out, neuron_2_add_20_out, neuron_2_add_21_out, neuron_2_add_22_out, neuron_2_add_23_out;
wire [25:0] neuron_2_add_24_out, neuron_2_add_25_out, neuron_2_add_26_out, neuron_2_add_27_out;

wire [25:0] neuron_3_add_0_out, neuron_3_add_1_out, neuron_3_add_2_out, neuron_3_add_3_out, neuron_3_add_4_out, neuron_3_add_5_out;
wire [25:0] neuron_3_add_6_out, neuron_3_add_7_out, neuron_3_add_8_out, neuron_3_add_9_out, neuron_3_add_10_out, neuron_3_add_11_out;
wire [25:0] neuron_3_add_12_out, neuron_3_add_13_out, neuron_3_add_14_out, neuron_3_add_15_out, neuron_3_add_16_out, neuron_3_add_17_out;
wire [25:0] neuron_3_add_18_out, neuron_3_add_19_out, neuron_3_add_20_out, neuron_3_add_21_out, neuron_3_add_22_out, neuron_3_add_23_out;
wire [25:0] neuron_3_add_24_out, neuron_3_add_25_out, neuron_3_add_26_out, neuron_3_add_27_out;

wire [25:0] neuron_4_add_0_out, neuron_4_add_1_out, neuron_4_add_2_out, neuron_4_add_3_out, neuron_4_add_4_out, neuron_4_add_5_out;
wire [25:0] neuron_4_add_6_out, neuron_4_add_7_out, neuron_4_add_8_out, neuron_4_add_9_out, neuron_4_add_10_out, neuron_4_add_11_out;
wire [25:0] neuron_4_add_12_out, neuron_4_add_13_out, neuron_4_add_14_out, neuron_4_add_15_out, neuron_4_add_16_out, neuron_4_add_17_out;
wire [25:0] neuron_4_add_18_out, neuron_4_add_19_out, neuron_4_add_20_out, neuron_4_add_21_out, neuron_4_add_22_out, neuron_4_add_23_out;
wire [25:0] neuron_4_add_24_out, neuron_4_add_25_out, neuron_4_add_26_out, neuron_4_add_27_out;

wire [25:0] neuron_5_add_0_out, neuron_5_add_1_out, neuron_5_add_2_out, neuron_5_add_3_out, neuron_5_add_4_out, neuron_5_add_5_out;
wire [25:0] neuron_5_add_6_out, neuron_5_add_7_out, neuron_5_add_8_out, neuron_5_add_9_out, neuron_5_add_10_out, neuron_5_add_11_out;
wire [25:0] neuron_5_add_12_out, neuron_5_add_13_out, neuron_5_add_14_out, neuron_5_add_15_out, neuron_5_add_16_out, neuron_5_add_17_out;
wire [25:0] neuron_5_add_18_out, neuron_5_add_19_out, neuron_5_add_20_out, neuron_5_add_21_out, neuron_5_add_22_out, neuron_5_add_23_out;
wire [25:0] neuron_5_add_24_out, neuron_5_add_25_out, neuron_5_add_26_out, neuron_5_add_27_out;

wire [25:0] neuron_6_add_0_out, neuron_6_add_1_out, neuron_6_add_2_out, neuron_6_add_3_out, neuron_6_add_4_out, neuron_6_add_5_out;
wire [25:0] neuron_6_add_6_out, neuron_6_add_7_out, neuron_6_add_8_out, neuron_6_add_9_out, neuron_6_add_10_out, neuron_6_add_11_out;
wire [25:0] neuron_6_add_12_out, neuron_6_add_13_out, neuron_6_add_14_out, neuron_6_add_15_out, neuron_6_add_16_out, neuron_6_add_17_out;
wire [25:0] neuron_6_add_18_out, neuron_6_add_19_out, neuron_6_add_20_out, neuron_6_add_21_out, neuron_6_add_22_out, neuron_6_add_23_out;
wire [25:0] neuron_6_add_24_out, neuron_6_add_25_out, neuron_6_add_26_out, neuron_6_add_27_out;

wire [25:0] neuron_7_add_0_out, neuron_7_add_1_out, neuron_7_add_2_out, neuron_7_add_3_out, neuron_7_add_4_out, neuron_7_add_5_out;
wire [25:0] neuron_7_add_6_out, neuron_7_add_7_out, neuron_7_add_8_out, neuron_7_add_9_out, neuron_7_add_10_out, neuron_7_add_11_out;
wire [25:0] neuron_7_add_12_out, neuron_7_add_13_out, neuron_7_add_14_out, neuron_7_add_15_out, neuron_7_add_16_out, neuron_7_add_17_out;
wire [25:0] neuron_7_add_18_out, neuron_7_add_19_out, neuron_7_add_20_out, neuron_7_add_21_out, neuron_7_add_22_out, neuron_7_add_23_out;
wire [25:0] neuron_7_add_24_out, neuron_7_add_25_out, neuron_7_add_26_out, neuron_7_add_27_out;

wire [25:0] neuron_8_add_0_out, neuron_8_add_1_out, neuron_8_add_2_out, neuron_8_add_3_out, neuron_8_add_4_out, neuron_8_add_5_out;
wire [25:0] neuron_8_add_6_out, neuron_8_add_7_out, neuron_8_add_8_out, neuron_8_add_9_out, neuron_8_add_10_out, neuron_8_add_11_out;
wire [25:0] neuron_8_add_12_out, neuron_8_add_13_out, neuron_8_add_14_out, neuron_8_add_15_out, neuron_8_add_16_out, neuron_8_add_17_out;
wire [25:0] neuron_8_add_18_out, neuron_8_add_19_out, neuron_8_add_20_out, neuron_8_add_21_out, neuron_8_add_22_out, neuron_8_add_23_out;
wire [25:0] neuron_8_add_24_out, neuron_8_add_25_out, neuron_8_add_26_out, neuron_8_add_27_out;

wire [25:0] neuron_9_add_0_out, neuron_9_add_1_out, neuron_9_add_2_out, neuron_9_add_3_out, neuron_9_add_4_out, neuron_9_add_5_out;
wire [25:0] neuron_9_add_6_out, neuron_9_add_7_out, neuron_9_add_8_out, neuron_9_add_9_out, neuron_9_add_10_out, neuron_9_add_11_out;
wire [25:0] neuron_9_add_12_out, neuron_9_add_13_out, neuron_9_add_14_out, neuron_9_add_15_out, neuron_9_add_16_out, neuron_9_add_17_out;
wire [25:0] neuron_9_add_18_out, neuron_9_add_19_out, neuron_9_add_20_out, neuron_9_add_21_out, neuron_9_add_22_out, neuron_9_add_23_out;
wire [25:0] neuron_9_add_24_out, neuron_9_add_25_out, neuron_9_add_26_out, neuron_9_add_27_out;

// Instantiate neuron multipliers
// neuron 0
FixedPointMultiplier neuron_0_mul_0(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_0_w), .PixelPort(neuron_mul_0_p), .Output_syn(neuron_0_mul_0_out));
FixedPointMultiplier neuron_0_mul_1(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_1_w), .PixelPort(neuron_mul_1_p), .Output_syn(neuron_0_mul_1_out));
FixedPointMultiplier neuron_0_mul_2(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_2_w), .PixelPort(neuron_mul_2_p), .Output_syn(neuron_0_mul_2_out));
FixedPointMultiplier neuron_0_mul_3(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_3_w), .PixelPort(neuron_mul_3_p), .Output_syn(neuron_0_mul_3_out));
FixedPointMultiplier neuron_0_mul_4(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_4_w), .PixelPort(neuron_mul_4_p), .Output_syn(neuron_0_mul_4_out));
FixedPointMultiplier neuron_0_mul_5(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_5_w), .PixelPort(neuron_mul_5_p), .Output_syn(neuron_0_mul_5_out));
FixedPointMultiplier neuron_0_mul_6(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_6_w), .PixelPort(neuron_mul_6_p), .Output_syn(neuron_0_mul_6_out));
FixedPointMultiplier neuron_0_mul_7(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_7_w), .PixelPort(neuron_mul_7_p), .Output_syn(neuron_0_mul_7_out));
FixedPointMultiplier neuron_0_mul_8(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_8_w), .PixelPort(neuron_mul_8_p), .Output_syn(neuron_0_mul_8_out));
FixedPointMultiplier neuron_0_mul_9(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_9_w), .PixelPort(neuron_mul_9_p), .Output_syn(neuron_0_mul_9_out));
FixedPointMultiplier neuron_0_mul_10(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_10_w), .PixelPort(neuron_mul_10_p), .Output_syn(neuron_0_mul_10_out));
FixedPointMultiplier neuron_0_mul_11(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_11_w), .PixelPort(neuron_mul_11_p), .Output_syn(neuron_0_mul_11_out));
FixedPointMultiplier neuron_0_mul_12(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_12_w), .PixelPort(neuron_mul_12_p), .Output_syn(neuron_0_mul_12_out));
FixedPointMultiplier neuron_0_mul_13(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_13_w), .PixelPort(neuron_mul_13_p), .Output_syn(neuron_0_mul_13_out));
FixedPointMultiplier neuron_0_mul_14(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_14_w), .PixelPort(neuron_mul_14_p), .Output_syn(neuron_0_mul_14_out));
FixedPointMultiplier neuron_0_mul_15(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_15_w), .PixelPort(neuron_mul_15_p), .Output_syn(neuron_0_mul_15_out));
FixedPointMultiplier neuron_0_mul_16(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_16_w), .PixelPort(neuron_mul_16_p), .Output_syn(neuron_0_mul_16_out));
FixedPointMultiplier neuron_0_mul_17(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_17_w), .PixelPort(neuron_mul_17_p), .Output_syn(neuron_0_mul_17_out));
FixedPointMultiplier neuron_0_mul_18(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_18_w), .PixelPort(neuron_mul_18_p), .Output_syn(neuron_0_mul_18_out));
FixedPointMultiplier neuron_0_mul_19(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_19_w), .PixelPort(neuron_mul_19_p), .Output_syn(neuron_0_mul_19_out));
FixedPointMultiplier neuron_0_mul_20(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_20_w), .PixelPort(neuron_mul_20_p), .Output_syn(neuron_0_mul_20_out));
FixedPointMultiplier neuron_0_mul_21(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_21_w), .PixelPort(neuron_mul_21_p), .Output_syn(neuron_0_mul_21_out));
FixedPointMultiplier neuron_0_mul_22(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_22_w), .PixelPort(neuron_mul_22_p), .Output_syn(neuron_0_mul_22_out));
FixedPointMultiplier neuron_0_mul_23(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_23_w), .PixelPort(neuron_mul_23_p), .Output_syn(neuron_0_mul_23_out));
FixedPointMultiplier neuron_0_mul_24(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_24_w), .PixelPort(neuron_mul_24_p), .Output_syn(neuron_0_mul_24_out));
FixedPointMultiplier neuron_0_mul_25(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_25_w), .PixelPort(neuron_mul_25_p), .Output_syn(neuron_0_mul_25_out));
FixedPointMultiplier neuron_0_mul_26(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_26_w), .PixelPort(neuron_mul_26_p), .Output_syn(neuron_0_mul_26_out));
FixedPointMultiplier neuron_0_mul_27(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_0_mul_27_w), .PixelPort(neuron_mul_27_p), .Output_syn(neuron_0_mul_27_out));

// neuron 1
FixedPointMultiplier neuron_1_mul_0(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_0_w), .PixelPort(neuron_mul_0_p), .Output_syn(neuron_1_mul_0_out));
FixedPointMultiplier neuron_1_mul_1(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_1_w), .PixelPort(neuron_mul_1_p), .Output_syn(neuron_1_mul_1_out));
FixedPointMultiplier neuron_1_mul_2(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_2_w), .PixelPort(neuron_mul_2_p), .Output_syn(neuron_1_mul_2_out));
FixedPointMultiplier neuron_1_mul_3(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_3_w), .PixelPort(neuron_mul_3_p), .Output_syn(neuron_1_mul_3_out));
FixedPointMultiplier neuron_1_mul_4(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_4_w), .PixelPort(neuron_mul_4_p), .Output_syn(neuron_1_mul_4_out));
FixedPointMultiplier neuron_1_mul_5(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_5_w), .PixelPort(neuron_mul_5_p), .Output_syn(neuron_1_mul_5_out));
FixedPointMultiplier neuron_1_mul_6(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_6_w), .PixelPort(neuron_mul_6_p), .Output_syn(neuron_1_mul_6_out));
FixedPointMultiplier neuron_1_mul_7(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_7_w), .PixelPort(neuron_mul_7_p), .Output_syn(neuron_1_mul_7_out));
FixedPointMultiplier neuron_1_mul_8(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_8_w), .PixelPort(neuron_mul_8_p), .Output_syn(neuron_1_mul_8_out));
FixedPointMultiplier neuron_1_mul_9(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_9_w), .PixelPort(neuron_mul_9_p), .Output_syn(neuron_1_mul_9_out));
FixedPointMultiplier neuron_1_mul_10(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_10_w), .PixelPort(neuron_mul_10_p), .Output_syn(neuron_1_mul_10_out));
FixedPointMultiplier neuron_1_mul_11(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_11_w), .PixelPort(neuron_mul_11_p), .Output_syn(neuron_1_mul_11_out));
FixedPointMultiplier neuron_1_mul_12(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_12_w), .PixelPort(neuron_mul_12_p), .Output_syn(neuron_1_mul_12_out));
FixedPointMultiplier neuron_1_mul_13(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_13_w), .PixelPort(neuron_mul_13_p), .Output_syn(neuron_1_mul_13_out));
FixedPointMultiplier neuron_1_mul_14(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_14_w), .PixelPort(neuron_mul_14_p), .Output_syn(neuron_1_mul_14_out));
FixedPointMultiplier neuron_1_mul_15(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_15_w), .PixelPort(neuron_mul_15_p), .Output_syn(neuron_1_mul_15_out));
FixedPointMultiplier neuron_1_mul_16(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_16_w), .PixelPort(neuron_mul_16_p), .Output_syn(neuron_1_mul_16_out));
FixedPointMultiplier neuron_1_mul_17(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_17_w), .PixelPort(neuron_mul_17_p), .Output_syn(neuron_1_mul_17_out));
FixedPointMultiplier neuron_1_mul_18(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_18_w), .PixelPort(neuron_mul_18_p), .Output_syn(neuron_1_mul_18_out));
FixedPointMultiplier neuron_1_mul_19(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_19_w), .PixelPort(neuron_mul_19_p), .Output_syn(neuron_1_mul_19_out));
FixedPointMultiplier neuron_1_mul_20(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_20_w), .PixelPort(neuron_mul_20_p), .Output_syn(neuron_1_mul_20_out));
FixedPointMultiplier neuron_1_mul_21(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_21_w), .PixelPort(neuron_mul_21_p), .Output_syn(neuron_1_mul_21_out));
FixedPointMultiplier neuron_1_mul_22(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_22_w), .PixelPort(neuron_mul_22_p), .Output_syn(neuron_1_mul_22_out));
FixedPointMultiplier neuron_1_mul_23(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_23_w), .PixelPort(neuron_mul_23_p), .Output_syn(neuron_1_mul_23_out));
FixedPointMultiplier neuron_1_mul_24(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_24_w), .PixelPort(neuron_mul_24_p), .Output_syn(neuron_1_mul_24_out));
FixedPointMultiplier neuron_1_mul_25(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_25_w), .PixelPort(neuron_mul_25_p), .Output_syn(neuron_1_mul_25_out));
FixedPointMultiplier neuron_1_mul_26(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_26_w), .PixelPort(neuron_mul_26_p), .Output_syn(neuron_1_mul_26_out));
FixedPointMultiplier neuron_1_mul_27(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_1_mul_27_w), .PixelPort(neuron_mul_27_p), .Output_syn(neuron_1_mul_27_out));

// neuron 2
FixedPointMultiplier neuron_2_mul_0(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_0_w), .PixelPort(neuron_mul_0_p), .Output_syn(neuron_2_mul_0_out));
FixedPointMultiplier neuron_2_mul_1(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_1_w), .PixelPort(neuron_mul_1_p), .Output_syn(neuron_2_mul_1_out));
FixedPointMultiplier neuron_2_mul_2(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_2_w), .PixelPort(neuron_mul_2_p), .Output_syn(neuron_2_mul_2_out));
FixedPointMultiplier neuron_2_mul_3(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_3_w), .PixelPort(neuron_mul_3_p), .Output_syn(neuron_2_mul_3_out));
FixedPointMultiplier neuron_2_mul_4(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_4_w), .PixelPort(neuron_mul_4_p), .Output_syn(neuron_2_mul_4_out));
FixedPointMultiplier neuron_2_mul_5(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_5_w), .PixelPort(neuron_mul_5_p), .Output_syn(neuron_2_mul_5_out));
FixedPointMultiplier neuron_2_mul_6(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_6_w), .PixelPort(neuron_mul_6_p), .Output_syn(neuron_2_mul_6_out));
FixedPointMultiplier neuron_2_mul_7(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_7_w), .PixelPort(neuron_mul_7_p), .Output_syn(neuron_2_mul_7_out));
FixedPointMultiplier neuron_2_mul_8(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_8_w), .PixelPort(neuron_mul_8_p), .Output_syn(neuron_2_mul_8_out));
FixedPointMultiplier neuron_2_mul_9(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_9_w), .PixelPort(neuron_mul_9_p), .Output_syn(neuron_2_mul_9_out));
FixedPointMultiplier neuron_2_mul_10(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_10_w), .PixelPort(neuron_mul_10_p), .Output_syn(neuron_2_mul_10_out));
FixedPointMultiplier neuron_2_mul_11(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_11_w), .PixelPort(neuron_mul_11_p), .Output_syn(neuron_2_mul_11_out));
FixedPointMultiplier neuron_2_mul_12(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_12_w), .PixelPort(neuron_mul_12_p), .Output_syn(neuron_2_mul_12_out));
FixedPointMultiplier neuron_2_mul_13(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_13_w), .PixelPort(neuron_mul_13_p), .Output_syn(neuron_2_mul_13_out));
FixedPointMultiplier neuron_2_mul_14(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_14_w), .PixelPort(neuron_mul_14_p), .Output_syn(neuron_2_mul_14_out));
FixedPointMultiplier neuron_2_mul_15(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_15_w), .PixelPort(neuron_mul_15_p), .Output_syn(neuron_2_mul_15_out));
FixedPointMultiplier neuron_2_mul_16(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_16_w), .PixelPort(neuron_mul_16_p), .Output_syn(neuron_2_mul_16_out));
FixedPointMultiplier neuron_2_mul_17(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_17_w), .PixelPort(neuron_mul_17_p), .Output_syn(neuron_2_mul_17_out));
FixedPointMultiplier neuron_2_mul_18(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_18_w), .PixelPort(neuron_mul_18_p), .Output_syn(neuron_2_mul_18_out));
FixedPointMultiplier neuron_2_mul_19(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_19_w), .PixelPort(neuron_mul_19_p), .Output_syn(neuron_2_mul_19_out));
FixedPointMultiplier neuron_2_mul_20(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_20_w), .PixelPort(neuron_mul_20_p), .Output_syn(neuron_2_mul_20_out));
FixedPointMultiplier neuron_2_mul_21(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_21_w), .PixelPort(neuron_mul_21_p), .Output_syn(neuron_2_mul_21_out));
FixedPointMultiplier neuron_2_mul_22(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_22_w), .PixelPort(neuron_mul_22_p), .Output_syn(neuron_2_mul_22_out));
FixedPointMultiplier neuron_2_mul_23(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_23_w), .PixelPort(neuron_mul_23_p), .Output_syn(neuron_2_mul_23_out));
FixedPointMultiplier neuron_2_mul_24(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_24_w), .PixelPort(neuron_mul_24_p), .Output_syn(neuron_2_mul_24_out));
FixedPointMultiplier neuron_2_mul_25(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_25_w), .PixelPort(neuron_mul_25_p), .Output_syn(neuron_2_mul_25_out));
FixedPointMultiplier neuron_2_mul_26(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_26_w), .PixelPort(neuron_mul_26_p), .Output_syn(neuron_2_mul_26_out));
FixedPointMultiplier neuron_2_mul_27(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_2_mul_27_w), .PixelPort(neuron_mul_27_p), .Output_syn(neuron_2_mul_27_out));

// neuron 3
FixedPointMultiplier neuron_3_mul_0(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_0_w), .PixelPort(neuron_mul_0_p), .Output_syn(neuron_3_mul_0_out));
FixedPointMultiplier neuron_3_mul_1(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_1_w), .PixelPort(neuron_mul_1_p), .Output_syn(neuron_3_mul_1_out));
FixedPointMultiplier neuron_3_mul_2(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_2_w), .PixelPort(neuron_mul_2_p), .Output_syn(neuron_3_mul_2_out));
FixedPointMultiplier neuron_3_mul_3(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_3_w), .PixelPort(neuron_mul_3_p), .Output_syn(neuron_3_mul_3_out));
FixedPointMultiplier neuron_3_mul_4(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_4_w), .PixelPort(neuron_mul_4_p), .Output_syn(neuron_3_mul_4_out));
FixedPointMultiplier neuron_3_mul_5(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_5_w), .PixelPort(neuron_mul_5_p), .Output_syn(neuron_3_mul_5_out));
FixedPointMultiplier neuron_3_mul_6(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_6_w), .PixelPort(neuron_mul_6_p), .Output_syn(neuron_3_mul_6_out));
FixedPointMultiplier neuron_3_mul_7(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_7_w), .PixelPort(neuron_mul_7_p), .Output_syn(neuron_3_mul_7_out));
FixedPointMultiplier neuron_3_mul_8(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_8_w), .PixelPort(neuron_mul_8_p), .Output_syn(neuron_3_mul_8_out));
FixedPointMultiplier neuron_3_mul_9(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_9_w), .PixelPort(neuron_mul_9_p), .Output_syn(neuron_3_mul_9_out));
FixedPointMultiplier neuron_3_mul_10(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_10_w), .PixelPort(neuron_mul_10_p), .Output_syn(neuron_3_mul_10_out));
FixedPointMultiplier neuron_3_mul_11(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_11_w), .PixelPort(neuron_mul_11_p), .Output_syn(neuron_3_mul_11_out));
FixedPointMultiplier neuron_3_mul_12(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_12_w), .PixelPort(neuron_mul_12_p), .Output_syn(neuron_3_mul_12_out));
FixedPointMultiplier neuron_3_mul_13(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_13_w), .PixelPort(neuron_mul_13_p), .Output_syn(neuron_3_mul_13_out));
FixedPointMultiplier neuron_3_mul_14(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_14_w), .PixelPort(neuron_mul_14_p), .Output_syn(neuron_3_mul_14_out));
FixedPointMultiplier neuron_3_mul_15(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_15_w), .PixelPort(neuron_mul_15_p), .Output_syn(neuron_3_mul_15_out));
FixedPointMultiplier neuron_3_mul_16(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_16_w), .PixelPort(neuron_mul_16_p), .Output_syn(neuron_3_mul_16_out));
FixedPointMultiplier neuron_3_mul_17(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_17_w), .PixelPort(neuron_mul_17_p), .Output_syn(neuron_3_mul_17_out));
FixedPointMultiplier neuron_3_mul_18(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_18_w), .PixelPort(neuron_mul_18_p), .Output_syn(neuron_3_mul_18_out));
FixedPointMultiplier neuron_3_mul_19(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_19_w), .PixelPort(neuron_mul_19_p), .Output_syn(neuron_3_mul_19_out));
FixedPointMultiplier neuron_3_mul_20(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_20_w), .PixelPort(neuron_mul_20_p), .Output_syn(neuron_3_mul_20_out));
FixedPointMultiplier neuron_3_mul_21(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_21_w), .PixelPort(neuron_mul_21_p), .Output_syn(neuron_3_mul_21_out));
FixedPointMultiplier neuron_3_mul_22(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_22_w), .PixelPort(neuron_mul_22_p), .Output_syn(neuron_3_mul_22_out));
FixedPointMultiplier neuron_3_mul_23(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_23_w), .PixelPort(neuron_mul_23_p), .Output_syn(neuron_3_mul_23_out));
FixedPointMultiplier neuron_3_mul_24(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_24_w), .PixelPort(neuron_mul_24_p), .Output_syn(neuron_3_mul_24_out));
FixedPointMultiplier neuron_3_mul_25(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_25_w), .PixelPort(neuron_mul_25_p), .Output_syn(neuron_3_mul_25_out));
FixedPointMultiplier neuron_3_mul_26(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_26_w), .PixelPort(neuron_mul_26_p), .Output_syn(neuron_3_mul_26_out));
FixedPointMultiplier neuron_3_mul_27(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_3_mul_27_w), .PixelPort(neuron_mul_27_p), .Output_syn(neuron_3_mul_27_out));

// neuron 4
FixedPointMultiplier neuron_4_mul_0(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_0_w), .PixelPort(neuron_mul_0_p), .Output_syn(neuron_4_mul_0_out));
FixedPointMultiplier neuron_4_mul_1(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_1_w), .PixelPort(neuron_mul_1_p), .Output_syn(neuron_4_mul_1_out));
FixedPointMultiplier neuron_4_mul_2(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_2_w), .PixelPort(neuron_mul_2_p), .Output_syn(neuron_4_mul_2_out));
FixedPointMultiplier neuron_4_mul_3(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_3_w), .PixelPort(neuron_mul_3_p), .Output_syn(neuron_4_mul_3_out));
FixedPointMultiplier neuron_4_mul_4(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_4_w), .PixelPort(neuron_mul_4_p), .Output_syn(neuron_4_mul_4_out));
FixedPointMultiplier neuron_4_mul_5(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_5_w), .PixelPort(neuron_mul_5_p), .Output_syn(neuron_4_mul_5_out));
FixedPointMultiplier neuron_4_mul_6(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_6_w), .PixelPort(neuron_mul_6_p), .Output_syn(neuron_4_mul_6_out));
FixedPointMultiplier neuron_4_mul_7(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_7_w), .PixelPort(neuron_mul_7_p), .Output_syn(neuron_4_mul_7_out));
FixedPointMultiplier neuron_4_mul_8(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_8_w), .PixelPort(neuron_mul_8_p), .Output_syn(neuron_4_mul_8_out));
FixedPointMultiplier neuron_4_mul_9(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_9_w), .PixelPort(neuron_mul_9_p), .Output_syn(neuron_4_mul_9_out));
FixedPointMultiplier neuron_4_mul_10(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_10_w), .PixelPort(neuron_mul_10_p), .Output_syn(neuron_4_mul_10_out));
FixedPointMultiplier neuron_4_mul_11(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_11_w), .PixelPort(neuron_mul_11_p), .Output_syn(neuron_4_mul_11_out));
FixedPointMultiplier neuron_4_mul_12(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_12_w), .PixelPort(neuron_mul_12_p), .Output_syn(neuron_4_mul_12_out));
FixedPointMultiplier neuron_4_mul_13(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_13_w), .PixelPort(neuron_mul_13_p), .Output_syn(neuron_4_mul_13_out));
FixedPointMultiplier neuron_4_mul_14(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_14_w), .PixelPort(neuron_mul_14_p), .Output_syn(neuron_4_mul_14_out));
FixedPointMultiplier neuron_4_mul_15(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_15_w), .PixelPort(neuron_mul_15_p), .Output_syn(neuron_4_mul_15_out));
FixedPointMultiplier neuron_4_mul_16(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_16_w), .PixelPort(neuron_mul_16_p), .Output_syn(neuron_4_mul_16_out));
FixedPointMultiplier neuron_4_mul_17(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_17_w), .PixelPort(neuron_mul_17_p), .Output_syn(neuron_4_mul_17_out));
FixedPointMultiplier neuron_4_mul_18(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_18_w), .PixelPort(neuron_mul_18_p), .Output_syn(neuron_4_mul_18_out));
FixedPointMultiplier neuron_4_mul_19(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_19_w), .PixelPort(neuron_mul_19_p), .Output_syn(neuron_4_mul_19_out));
FixedPointMultiplier neuron_4_mul_20(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_20_w), .PixelPort(neuron_mul_20_p), .Output_syn(neuron_4_mul_20_out));
FixedPointMultiplier neuron_4_mul_21(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_21_w), .PixelPort(neuron_mul_21_p), .Output_syn(neuron_4_mul_21_out));
FixedPointMultiplier neuron_4_mul_22(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_22_w), .PixelPort(neuron_mul_22_p), .Output_syn(neuron_4_mul_22_out));
FixedPointMultiplier neuron_4_mul_23(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_23_w), .PixelPort(neuron_mul_23_p), .Output_syn(neuron_4_mul_23_out));
FixedPointMultiplier neuron_4_mul_24(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_24_w), .PixelPort(neuron_mul_24_p), .Output_syn(neuron_4_mul_24_out));
FixedPointMultiplier neuron_4_mul_25(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_25_w), .PixelPort(neuron_mul_25_p), .Output_syn(neuron_4_mul_25_out));
FixedPointMultiplier neuron_4_mul_26(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_26_w), .PixelPort(neuron_mul_26_p), .Output_syn(neuron_4_mul_26_out));
FixedPointMultiplier neuron_4_mul_27(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_4_mul_27_w), .PixelPort(neuron_mul_27_p), .Output_syn(neuron_4_mul_27_out));

// neuron 5
FixedPointMultiplier neuron_5_mul_0(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_0_w), .PixelPort(neuron_mul_0_p), .Output_syn(neuron_5_mul_0_out));
FixedPointMultiplier neuron_5_mul_1(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_1_w), .PixelPort(neuron_mul_1_p), .Output_syn(neuron_5_mul_1_out));
FixedPointMultiplier neuron_5_mul_2(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_2_w), .PixelPort(neuron_mul_2_p), .Output_syn(neuron_5_mul_2_out));
FixedPointMultiplier neuron_5_mul_3(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_3_w), .PixelPort(neuron_mul_3_p), .Output_syn(neuron_5_mul_3_out));
FixedPointMultiplier neuron_5_mul_4(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_4_w), .PixelPort(neuron_mul_4_p), .Output_syn(neuron_5_mul_4_out));
FixedPointMultiplier neuron_5_mul_5(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_5_w), .PixelPort(neuron_mul_5_p), .Output_syn(neuron_5_mul_5_out));
FixedPointMultiplier neuron_5_mul_6(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_6_w), .PixelPort(neuron_mul_6_p), .Output_syn(neuron_5_mul_6_out));
FixedPointMultiplier neuron_5_mul_7(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_7_w), .PixelPort(neuron_mul_7_p), .Output_syn(neuron_5_mul_7_out));
FixedPointMultiplier neuron_5_mul_8(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_8_w), .PixelPort(neuron_mul_8_p), .Output_syn(neuron_5_mul_8_out));
FixedPointMultiplier neuron_5_mul_9(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_9_w), .PixelPort(neuron_mul_9_p), .Output_syn(neuron_5_mul_9_out));
FixedPointMultiplier neuron_5_mul_10(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_10_w), .PixelPort(neuron_mul_10_p), .Output_syn(neuron_5_mul_10_out));
FixedPointMultiplier neuron_5_mul_11(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_11_w), .PixelPort(neuron_mul_11_p), .Output_syn(neuron_5_mul_11_out));
FixedPointMultiplier neuron_5_mul_12(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_12_w), .PixelPort(neuron_mul_12_p), .Output_syn(neuron_5_mul_12_out));
FixedPointMultiplier neuron_5_mul_13(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_13_w), .PixelPort(neuron_mul_13_p), .Output_syn(neuron_5_mul_13_out));
FixedPointMultiplier neuron_5_mul_14(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_14_w), .PixelPort(neuron_mul_14_p), .Output_syn(neuron_5_mul_14_out));
FixedPointMultiplier neuron_5_mul_15(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_15_w), .PixelPort(neuron_mul_15_p), .Output_syn(neuron_5_mul_15_out));
FixedPointMultiplier neuron_5_mul_16(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_16_w), .PixelPort(neuron_mul_16_p), .Output_syn(neuron_5_mul_16_out));
FixedPointMultiplier neuron_5_mul_17(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_17_w), .PixelPort(neuron_mul_17_p), .Output_syn(neuron_5_mul_17_out));
FixedPointMultiplier neuron_5_mul_18(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_18_w), .PixelPort(neuron_mul_18_p), .Output_syn(neuron_5_mul_18_out));
FixedPointMultiplier neuron_5_mul_19(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_19_w), .PixelPort(neuron_mul_19_p), .Output_syn(neuron_5_mul_19_out));
FixedPointMultiplier neuron_5_mul_20(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_20_w), .PixelPort(neuron_mul_20_p), .Output_syn(neuron_5_mul_20_out));
FixedPointMultiplier neuron_5_mul_21(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_21_w), .PixelPort(neuron_mul_21_p), .Output_syn(neuron_5_mul_21_out));
FixedPointMultiplier neuron_5_mul_22(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_22_w), .PixelPort(neuron_mul_22_p), .Output_syn(neuron_5_mul_22_out));
FixedPointMultiplier neuron_5_mul_23(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_23_w), .PixelPort(neuron_mul_23_p), .Output_syn(neuron_5_mul_23_out));
FixedPointMultiplier neuron_5_mul_24(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_24_w), .PixelPort(neuron_mul_24_p), .Output_syn(neuron_5_mul_24_out));
FixedPointMultiplier neuron_5_mul_25(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_25_w), .PixelPort(neuron_mul_25_p), .Output_syn(neuron_5_mul_25_out));
FixedPointMultiplier neuron_5_mul_26(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_26_w), .PixelPort(neuron_mul_26_p), .Output_syn(neuron_5_mul_26_out));
FixedPointMultiplier neuron_5_mul_27(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_5_mul_27_w), .PixelPort(neuron_mul_27_p), .Output_syn(neuron_5_mul_27_out));

// neuron 6
FixedPointMultiplier neuron_6_mul_0(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_0_w), .PixelPort(neuron_mul_0_p), .Output_syn(neuron_6_mul_0_out));
FixedPointMultiplier neuron_6_mul_1(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_1_w), .PixelPort(neuron_mul_1_p), .Output_syn(neuron_6_mul_1_out));
FixedPointMultiplier neuron_6_mul_2(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_2_w), .PixelPort(neuron_mul_2_p), .Output_syn(neuron_6_mul_2_out));
FixedPointMultiplier neuron_6_mul_3(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_3_w), .PixelPort(neuron_mul_3_p), .Output_syn(neuron_6_mul_3_out));
FixedPointMultiplier neuron_6_mul_4(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_4_w), .PixelPort(neuron_mul_4_p), .Output_syn(neuron_6_mul_4_out));
FixedPointMultiplier neuron_6_mul_5(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_5_w), .PixelPort(neuron_mul_5_p), .Output_syn(neuron_6_mul_5_out));
FixedPointMultiplier neuron_6_mul_6(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_6_w), .PixelPort(neuron_mul_6_p), .Output_syn(neuron_6_mul_6_out));
FixedPointMultiplier neuron_6_mul_7(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_7_w), .PixelPort(neuron_mul_7_p), .Output_syn(neuron_6_mul_7_out));
FixedPointMultiplier neuron_6_mul_8(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_8_w), .PixelPort(neuron_mul_8_p), .Output_syn(neuron_6_mul_8_out));
FixedPointMultiplier neuron_6_mul_9(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_9_w), .PixelPort(neuron_mul_9_p), .Output_syn(neuron_6_mul_9_out));
FixedPointMultiplier neuron_6_mul_10(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_10_w), .PixelPort(neuron_mul_10_p), .Output_syn(neuron_6_mul_10_out));
FixedPointMultiplier neuron_6_mul_11(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_11_w), .PixelPort(neuron_mul_11_p), .Output_syn(neuron_6_mul_11_out));
FixedPointMultiplier neuron_6_mul_12(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_12_w), .PixelPort(neuron_mul_12_p), .Output_syn(neuron_6_mul_12_out));
FixedPointMultiplier neuron_6_mul_13(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_13_w), .PixelPort(neuron_mul_13_p), .Output_syn(neuron_6_mul_13_out));
FixedPointMultiplier neuron_6_mul_14(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_14_w), .PixelPort(neuron_mul_14_p), .Output_syn(neuron_6_mul_14_out));
FixedPointMultiplier neuron_6_mul_15(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_15_w), .PixelPort(neuron_mul_15_p), .Output_syn(neuron_6_mul_15_out));
FixedPointMultiplier neuron_6_mul_16(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_16_w), .PixelPort(neuron_mul_16_p), .Output_syn(neuron_6_mul_16_out));
FixedPointMultiplier neuron_6_mul_17(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_17_w), .PixelPort(neuron_mul_17_p), .Output_syn(neuron_6_mul_17_out));
FixedPointMultiplier neuron_6_mul_18(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_18_w), .PixelPort(neuron_mul_18_p), .Output_syn(neuron_6_mul_18_out));
FixedPointMultiplier neuron_6_mul_19(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_19_w), .PixelPort(neuron_mul_19_p), .Output_syn(neuron_6_mul_19_out));
FixedPointMultiplier neuron_6_mul_20(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_20_w), .PixelPort(neuron_mul_20_p), .Output_syn(neuron_6_mul_20_out));
FixedPointMultiplier neuron_6_mul_21(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_21_w), .PixelPort(neuron_mul_21_p), .Output_syn(neuron_6_mul_21_out));
FixedPointMultiplier neuron_6_mul_22(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_22_w), .PixelPort(neuron_mul_22_p), .Output_syn(neuron_6_mul_22_out));
FixedPointMultiplier neuron_6_mul_23(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_23_w), .PixelPort(neuron_mul_23_p), .Output_syn(neuron_6_mul_23_out));
FixedPointMultiplier neuron_6_mul_24(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_24_w), .PixelPort(neuron_mul_24_p), .Output_syn(neuron_6_mul_24_out));
FixedPointMultiplier neuron_6_mul_25(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_25_w), .PixelPort(neuron_mul_25_p), .Output_syn(neuron_6_mul_25_out));
FixedPointMultiplier neuron_6_mul_26(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_26_w), .PixelPort(neuron_mul_26_p), .Output_syn(neuron_6_mul_26_out));
FixedPointMultiplier neuron_6_mul_27(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_6_mul_27_w), .PixelPort(neuron_mul_27_p), .Output_syn(neuron_6_mul_27_out));

// neuron 7
FixedPointMultiplier neuron_7_mul_0(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_0_w), .PixelPort(neuron_mul_0_p), .Output_syn(neuron_7_mul_0_out));
FixedPointMultiplier neuron_7_mul_1(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_1_w), .PixelPort(neuron_mul_1_p), .Output_syn(neuron_7_mul_1_out));
FixedPointMultiplier neuron_7_mul_2(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_2_w), .PixelPort(neuron_mul_2_p), .Output_syn(neuron_7_mul_2_out));
FixedPointMultiplier neuron_7_mul_3(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_3_w), .PixelPort(neuron_mul_3_p), .Output_syn(neuron_7_mul_3_out));
FixedPointMultiplier neuron_7_mul_4(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_4_w), .PixelPort(neuron_mul_4_p), .Output_syn(neuron_7_mul_4_out));
FixedPointMultiplier neuron_7_mul_5(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_5_w), .PixelPort(neuron_mul_5_p), .Output_syn(neuron_7_mul_5_out));
FixedPointMultiplier neuron_7_mul_6(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_6_w), .PixelPort(neuron_mul_6_p), .Output_syn(neuron_7_mul_6_out));
FixedPointMultiplier neuron_7_mul_7(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_7_w), .PixelPort(neuron_mul_7_p), .Output_syn(neuron_7_mul_7_out));
FixedPointMultiplier neuron_7_mul_8(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_8_w), .PixelPort(neuron_mul_8_p), .Output_syn(neuron_7_mul_8_out));
FixedPointMultiplier neuron_7_mul_9(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_9_w), .PixelPort(neuron_mul_9_p), .Output_syn(neuron_7_mul_9_out));
FixedPointMultiplier neuron_7_mul_10(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_10_w), .PixelPort(neuron_mul_10_p), .Output_syn(neuron_7_mul_10_out));
FixedPointMultiplier neuron_7_mul_11(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_11_w), .PixelPort(neuron_mul_11_p), .Output_syn(neuron_7_mul_11_out));
FixedPointMultiplier neuron_7_mul_12(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_12_w), .PixelPort(neuron_mul_12_p), .Output_syn(neuron_7_mul_12_out));
FixedPointMultiplier neuron_7_mul_13(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_13_w), .PixelPort(neuron_mul_13_p), .Output_syn(neuron_7_mul_13_out));
FixedPointMultiplier neuron_7_mul_14(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_14_w), .PixelPort(neuron_mul_14_p), .Output_syn(neuron_7_mul_14_out));
FixedPointMultiplier neuron_7_mul_15(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_15_w), .PixelPort(neuron_mul_15_p), .Output_syn(neuron_7_mul_15_out));
FixedPointMultiplier neuron_7_mul_16(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_16_w), .PixelPort(neuron_mul_16_p), .Output_syn(neuron_7_mul_16_out));
FixedPointMultiplier neuron_7_mul_17(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_17_w), .PixelPort(neuron_mul_17_p), .Output_syn(neuron_7_mul_17_out));
FixedPointMultiplier neuron_7_mul_18(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_18_w), .PixelPort(neuron_mul_18_p), .Output_syn(neuron_7_mul_18_out));
FixedPointMultiplier neuron_7_mul_19(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_19_w), .PixelPort(neuron_mul_19_p), .Output_syn(neuron_7_mul_19_out));
FixedPointMultiplier neuron_7_mul_20(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_20_w), .PixelPort(neuron_mul_20_p), .Output_syn(neuron_7_mul_20_out));
FixedPointMultiplier neuron_7_mul_21(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_21_w), .PixelPort(neuron_mul_21_p), .Output_syn(neuron_7_mul_21_out));
FixedPointMultiplier neuron_7_mul_22(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_22_w), .PixelPort(neuron_mul_22_p), .Output_syn(neuron_7_mul_22_out));
FixedPointMultiplier neuron_7_mul_23(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_23_w), .PixelPort(neuron_mul_23_p), .Output_syn(neuron_7_mul_23_out));
FixedPointMultiplier neuron_7_mul_24(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_24_w), .PixelPort(neuron_mul_24_p), .Output_syn(neuron_7_mul_24_out));
FixedPointMultiplier neuron_7_mul_25(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_25_w), .PixelPort(neuron_mul_25_p), .Output_syn(neuron_7_mul_25_out));
FixedPointMultiplier neuron_7_mul_26(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_26_w), .PixelPort(neuron_mul_26_p), .Output_syn(neuron_7_mul_26_out));
FixedPointMultiplier neuron_7_mul_27(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_7_mul_27_w), .PixelPort(neuron_mul_27_p), .Output_syn(neuron_7_mul_27_out));

// neuron 8
FixedPointMultiplier neuron_8_mul_0(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_0_w), .PixelPort(neuron_mul_0_p), .Output_syn(neuron_8_mul_0_out));
FixedPointMultiplier neuron_8_mul_1(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_1_w), .PixelPort(neuron_mul_1_p), .Output_syn(neuron_8_mul_1_out));
FixedPointMultiplier neuron_8_mul_2(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_2_w), .PixelPort(neuron_mul_2_p), .Output_syn(neuron_8_mul_2_out));
FixedPointMultiplier neuron_8_mul_3(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_3_w), .PixelPort(neuron_mul_3_p), .Output_syn(neuron_8_mul_3_out));
FixedPointMultiplier neuron_8_mul_4(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_4_w), .PixelPort(neuron_mul_4_p), .Output_syn(neuron_8_mul_4_out));
FixedPointMultiplier neuron_8_mul_5(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_5_w), .PixelPort(neuron_mul_5_p), .Output_syn(neuron_8_mul_5_out));
FixedPointMultiplier neuron_8_mul_6(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_6_w), .PixelPort(neuron_mul_6_p), .Output_syn(neuron_8_mul_6_out));
FixedPointMultiplier neuron_8_mul_7(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_7_w), .PixelPort(neuron_mul_7_p), .Output_syn(neuron_8_mul_7_out));
FixedPointMultiplier neuron_8_mul_8(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_8_w), .PixelPort(neuron_mul_8_p), .Output_syn(neuron_8_mul_8_out));
FixedPointMultiplier neuron_8_mul_9(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_9_w), .PixelPort(neuron_mul_9_p), .Output_syn(neuron_8_mul_9_out));
FixedPointMultiplier neuron_8_mul_10(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_10_w), .PixelPort(neuron_mul_10_p), .Output_syn(neuron_8_mul_10_out));
FixedPointMultiplier neuron_8_mul_11(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_11_w), .PixelPort(neuron_mul_11_p), .Output_syn(neuron_8_mul_11_out));
FixedPointMultiplier neuron_8_mul_12(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_12_w), .PixelPort(neuron_mul_12_p), .Output_syn(neuron_8_mul_12_out));
FixedPointMultiplier neuron_8_mul_13(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_13_w), .PixelPort(neuron_mul_13_p), .Output_syn(neuron_8_mul_13_out));
FixedPointMultiplier neuron_8_mul_14(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_14_w), .PixelPort(neuron_mul_14_p), .Output_syn(neuron_8_mul_14_out));
FixedPointMultiplier neuron_8_mul_15(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_15_w), .PixelPort(neuron_mul_15_p), .Output_syn(neuron_8_mul_15_out));
FixedPointMultiplier neuron_8_mul_16(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_16_w), .PixelPort(neuron_mul_16_p), .Output_syn(neuron_8_mul_16_out));
FixedPointMultiplier neuron_8_mul_17(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_17_w), .PixelPort(neuron_mul_17_p), .Output_syn(neuron_8_mul_17_out));
FixedPointMultiplier neuron_8_mul_18(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_18_w), .PixelPort(neuron_mul_18_p), .Output_syn(neuron_8_mul_18_out));
FixedPointMultiplier neuron_8_mul_19(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_19_w), .PixelPort(neuron_mul_19_p), .Output_syn(neuron_8_mul_19_out));
FixedPointMultiplier neuron_8_mul_20(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_20_w), .PixelPort(neuron_mul_20_p), .Output_syn(neuron_8_mul_20_out));
FixedPointMultiplier neuron_8_mul_21(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_21_w), .PixelPort(neuron_mul_21_p), .Output_syn(neuron_8_mul_21_out));
FixedPointMultiplier neuron_8_mul_22(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_22_w), .PixelPort(neuron_mul_22_p), .Output_syn(neuron_8_mul_22_out));
FixedPointMultiplier neuron_8_mul_23(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_23_w), .PixelPort(neuron_mul_23_p), .Output_syn(neuron_8_mul_23_out));
FixedPointMultiplier neuron_8_mul_24(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_24_w), .PixelPort(neuron_mul_24_p), .Output_syn(neuron_8_mul_24_out));
FixedPointMultiplier neuron_8_mul_25(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_25_w), .PixelPort(neuron_mul_25_p), .Output_syn(neuron_8_mul_25_out));
FixedPointMultiplier neuron_8_mul_26(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_26_w), .PixelPort(neuron_mul_26_p), .Output_syn(neuron_8_mul_26_out));
FixedPointMultiplier neuron_8_mul_27(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_8_mul_27_w), .PixelPort(neuron_mul_27_p), .Output_syn(neuron_8_mul_27_out));

// neuron 9
FixedPointMultiplier neuron_9_mul_0(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_0_w), .PixelPort(neuron_mul_0_p), .Output_syn(neuron_9_mul_0_out));
FixedPointMultiplier neuron_9_mul_1(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_1_w), .PixelPort(neuron_mul_1_p), .Output_syn(neuron_9_mul_1_out));
FixedPointMultiplier neuron_9_mul_2(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_2_w), .PixelPort(neuron_mul_2_p), .Output_syn(neuron_9_mul_2_out));
FixedPointMultiplier neuron_9_mul_3(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_3_w), .PixelPort(neuron_mul_3_p), .Output_syn(neuron_9_mul_3_out));
FixedPointMultiplier neuron_9_mul_4(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_4_w), .PixelPort(neuron_mul_4_p), .Output_syn(neuron_9_mul_4_out));
FixedPointMultiplier neuron_9_mul_5(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_5_w), .PixelPort(neuron_mul_5_p), .Output_syn(neuron_9_mul_5_out));
FixedPointMultiplier neuron_9_mul_6(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_6_w), .PixelPort(neuron_mul_6_p), .Output_syn(neuron_9_mul_6_out));
FixedPointMultiplier neuron_9_mul_7(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_7_w), .PixelPort(neuron_mul_7_p), .Output_syn(neuron_9_mul_7_out));
FixedPointMultiplier neuron_9_mul_8(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_8_w), .PixelPort(neuron_mul_8_p), .Output_syn(neuron_9_mul_8_out));
FixedPointMultiplier neuron_9_mul_9(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_9_w), .PixelPort(neuron_mul_9_p), .Output_syn(neuron_9_mul_9_out));
FixedPointMultiplier neuron_9_mul_10(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_10_w), .PixelPort(neuron_mul_10_p), .Output_syn(neuron_9_mul_10_out));
FixedPointMultiplier neuron_9_mul_11(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_11_w), .PixelPort(neuron_mul_11_p), .Output_syn(neuron_9_mul_11_out));
FixedPointMultiplier neuron_9_mul_12(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_12_w), .PixelPort(neuron_mul_12_p), .Output_syn(neuron_9_mul_12_out));
FixedPointMultiplier neuron_9_mul_13(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_13_w), .PixelPort(neuron_mul_13_p), .Output_syn(neuron_9_mul_13_out));
FixedPointMultiplier neuron_9_mul_14(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_14_w), .PixelPort(neuron_mul_14_p), .Output_syn(neuron_9_mul_14_out));
FixedPointMultiplier neuron_9_mul_15(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_15_w), .PixelPort(neuron_mul_15_p), .Output_syn(neuron_9_mul_15_out));
FixedPointMultiplier neuron_9_mul_16(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_16_w), .PixelPort(neuron_mul_16_p), .Output_syn(neuron_9_mul_16_out));
FixedPointMultiplier neuron_9_mul_17(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_17_w), .PixelPort(neuron_mul_17_p), .Output_syn(neuron_9_mul_17_out));
FixedPointMultiplier neuron_9_mul_18(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_18_w), .PixelPort(neuron_mul_18_p), .Output_syn(neuron_9_mul_18_out));
FixedPointMultiplier neuron_9_mul_19(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_19_w), .PixelPort(neuron_mul_19_p), .Output_syn(neuron_9_mul_19_out));
FixedPointMultiplier neuron_9_mul_20(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_20_w), .PixelPort(neuron_mul_20_p), .Output_syn(neuron_9_mul_20_out));
FixedPointMultiplier neuron_9_mul_21(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_21_w), .PixelPort(neuron_mul_21_p), .Output_syn(neuron_9_mul_21_out));
FixedPointMultiplier neuron_9_mul_22(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_22_w), .PixelPort(neuron_mul_22_p), .Output_syn(neuron_9_mul_22_out));
FixedPointMultiplier neuron_9_mul_23(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_23_w), .PixelPort(neuron_mul_23_p), .Output_syn(neuron_9_mul_23_out));
FixedPointMultiplier neuron_9_mul_24(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_24_w), .PixelPort(neuron_mul_24_p), .Output_syn(neuron_9_mul_24_out));
FixedPointMultiplier neuron_9_mul_25(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_25_w), .PixelPort(neuron_mul_25_p), .Output_syn(neuron_9_mul_25_out));
FixedPointMultiplier neuron_9_mul_26(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_26_w), .PixelPort(neuron_mul_26_p), .Output_syn(neuron_9_mul_26_out));
FixedPointMultiplier neuron_9_mul_27(.clk(neuron_clk), .GlobalReset(globalreset), .WeightPort(neuron_9_mul_27_w), .PixelPort(neuron_mul_27_p), .Output_syn(neuron_9_mul_27_out));

// Instantiate neuron adders
// neuron 0
FixedPointAdder neuron_0_add_0(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_0_p1), .Port2(neuron_0_add_0_p2), .Output_syn(neuron_0_add_0_out));
FixedPointAdder neuron_0_add_1(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_1_p1), .Port2(neuron_0_add_1_p2), .Output_syn(neuron_0_add_1_out));
FixedPointAdder neuron_0_add_2(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_2_p1), .Port2(neuron_0_add_2_p2), .Output_syn(neuron_0_add_2_out));
FixedPointAdder neuron_0_add_3(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_3_p1), .Port2(neuron_0_add_3_p2), .Output_syn(neuron_0_add_3_out));
FixedPointAdder neuron_0_add_4(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_4_p1), .Port2(neuron_0_add_4_p2), .Output_syn(neuron_0_add_4_out));
FixedPointAdder neuron_0_add_5(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_5_p1), .Port2(neuron_0_add_5_p2), .Output_syn(neuron_0_add_5_out));
FixedPointAdder neuron_0_add_6(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_6_p1), .Port2(neuron_0_add_6_p2), .Output_syn(neuron_0_add_6_out));
FixedPointAdder neuron_0_add_7(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_7_p1), .Port2(neuron_0_add_7_p2), .Output_syn(neuron_0_add_7_out));
FixedPointAdder neuron_0_add_8(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_8_p1), .Port2(neuron_0_add_8_p2), .Output_syn(neuron_0_add_8_out));
FixedPointAdder neuron_0_add_9(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_9_p1), .Port2(neuron_0_add_9_p2), .Output_syn(neuron_0_add_9_out));
FixedPointAdder neuron_0_add_10(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_10_p1), .Port2(neuron_0_add_10_p2), .Output_syn(neuron_0_add_10_out));
FixedPointAdder neuron_0_add_11(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_11_p1), .Port2(neuron_0_add_11_p2), .Output_syn(neuron_0_add_11_out));
FixedPointAdder neuron_0_add_12(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_12_p1), .Port2(neuron_0_add_12_p2), .Output_syn(neuron_0_add_12_out));
FixedPointAdder neuron_0_add_13(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_13_p1), .Port2(neuron_0_add_13_p2), .Output_syn(neuron_0_add_13_out));
FixedPointAdder neuron_0_add_14(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_14_p1), .Port2(neuron_0_add_14_p2), .Output_syn(neuron_0_add_14_out));
FixedPointAdder neuron_0_add_15(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_15_p1), .Port2(neuron_0_add_15_p2), .Output_syn(neuron_0_add_15_out));
FixedPointAdder neuron_0_add_16(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_16_p1), .Port2(neuron_0_add_16_p2), .Output_syn(neuron_0_add_16_out));
FixedPointAdder neuron_0_add_17(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_17_p1), .Port2(neuron_0_add_17_p2), .Output_syn(neuron_0_add_17_out));
FixedPointAdder neuron_0_add_18(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_18_p1), .Port2(neuron_0_add_18_p2), .Output_syn(neuron_0_add_18_out));
FixedPointAdder neuron_0_add_19(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_19_p1), .Port2(neuron_0_add_19_p2), .Output_syn(neuron_0_add_19_out));
FixedPointAdder neuron_0_add_20(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_20_p1), .Port2(neuron_0_add_20_p2), .Output_syn(neuron_0_add_20_out));
FixedPointAdder neuron_0_add_21(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_21_p1), .Port2(neuron_0_add_21_p2), .Output_syn(neuron_0_add_21_out));
FixedPointAdder neuron_0_add_22(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_22_p1), .Port2(neuron_0_add_22_p2), .Output_syn(neuron_0_add_22_out));
FixedPointAdder neuron_0_add_23(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_23_p1), .Port2(neuron_0_add_23_p2), .Output_syn(neuron_0_add_23_out));
FixedPointAdder neuron_0_add_24(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_24_p1), .Port2(neuron_0_add_24_p2), .Output_syn(neuron_0_add_24_out));
FixedPointAdder neuron_0_add_25(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_25_p1), .Port2(neuron_0_add_25_p2), .Output_syn(neuron_0_add_25_out));
FixedPointAdder neuron_0_add_26(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_26_p1), .Port2(neuron_0_add_26_p2), .Output_syn(neuron_0_add_26_out));
FixedPointAdder neuron_0_add_27(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_0_add_27_p1), .Port2(neuron_0_add_27_p2), .Output_syn(neuron_0_add_27_out));

// neuron 1
FixedPointAdder neuron_1_add_0(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_0_p1), .Port2(neuron_1_add_0_p2), .Output_syn(neuron_1_add_0_out));
FixedPointAdder neuron_1_add_1(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_1_p1), .Port2(neuron_1_add_1_p2), .Output_syn(neuron_1_add_1_out));
FixedPointAdder neuron_1_add_2(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_2_p1), .Port2(neuron_1_add_2_p2), .Output_syn(neuron_1_add_2_out));
FixedPointAdder neuron_1_add_3(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_3_p1), .Port2(neuron_1_add_3_p2), .Output_syn(neuron_1_add_3_out));
FixedPointAdder neuron_1_add_4(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_4_p1), .Port2(neuron_1_add_4_p2), .Output_syn(neuron_1_add_4_out));
FixedPointAdder neuron_1_add_5(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_5_p1), .Port2(neuron_1_add_5_p2), .Output_syn(neuron_1_add_5_out));
FixedPointAdder neuron_1_add_6(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_6_p1), .Port2(neuron_1_add_6_p2), .Output_syn(neuron_1_add_6_out));
FixedPointAdder neuron_1_add_7(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_7_p1), .Port2(neuron_1_add_7_p2), .Output_syn(neuron_1_add_7_out));
FixedPointAdder neuron_1_add_8(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_8_p1), .Port2(neuron_1_add_8_p2), .Output_syn(neuron_1_add_8_out));
FixedPointAdder neuron_1_add_9(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_9_p1), .Port2(neuron_1_add_9_p2), .Output_syn(neuron_1_add_9_out));
FixedPointAdder neuron_1_add_10(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_10_p1), .Port2(neuron_1_add_10_p2), .Output_syn(neuron_1_add_10_out));
FixedPointAdder neuron_1_add_11(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_11_p1), .Port2(neuron_1_add_11_p2), .Output_syn(neuron_1_add_11_out));
FixedPointAdder neuron_1_add_12(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_12_p1), .Port2(neuron_1_add_12_p2), .Output_syn(neuron_1_add_12_out));
FixedPointAdder neuron_1_add_13(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_13_p1), .Port2(neuron_1_add_13_p2), .Output_syn(neuron_1_add_13_out));
FixedPointAdder neuron_1_add_14(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_14_p1), .Port2(neuron_1_add_14_p2), .Output_syn(neuron_1_add_14_out));
FixedPointAdder neuron_1_add_15(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_15_p1), .Port2(neuron_1_add_15_p2), .Output_syn(neuron_1_add_15_out));
FixedPointAdder neuron_1_add_16(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_16_p1), .Port2(neuron_1_add_16_p2), .Output_syn(neuron_1_add_16_out));
FixedPointAdder neuron_1_add_17(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_17_p1), .Port2(neuron_1_add_17_p2), .Output_syn(neuron_1_add_17_out));
FixedPointAdder neuron_1_add_18(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_18_p1), .Port2(neuron_1_add_18_p2), .Output_syn(neuron_1_add_18_out));
FixedPointAdder neuron_1_add_19(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_19_p1), .Port2(neuron_1_add_19_p2), .Output_syn(neuron_1_add_19_out));
FixedPointAdder neuron_1_add_20(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_20_p1), .Port2(neuron_1_add_20_p2), .Output_syn(neuron_1_add_20_out));
FixedPointAdder neuron_1_add_21(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_21_p1), .Port2(neuron_1_add_21_p2), .Output_syn(neuron_1_add_21_out));
FixedPointAdder neuron_1_add_22(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_22_p1), .Port2(neuron_1_add_22_p2), .Output_syn(neuron_1_add_22_out));
FixedPointAdder neuron_1_add_23(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_23_p1), .Port2(neuron_1_add_23_p2), .Output_syn(neuron_1_add_23_out));
FixedPointAdder neuron_1_add_24(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_24_p1), .Port2(neuron_1_add_24_p2), .Output_syn(neuron_1_add_24_out));
FixedPointAdder neuron_1_add_25(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_25_p1), .Port2(neuron_1_add_25_p2), .Output_syn(neuron_1_add_25_out));
FixedPointAdder neuron_1_add_26(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_26_p1), .Port2(neuron_1_add_26_p2), .Output_syn(neuron_1_add_26_out));
FixedPointAdder neuron_1_add_27(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_1_add_27_p1), .Port2(neuron_1_add_27_p2), .Output_syn(neuron_1_add_27_out));

// neuron 2
FixedPointAdder neuron_2_add_0(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_0_p1), .Port2(neuron_2_add_0_p2), .Output_syn(neuron_2_add_0_out));
FixedPointAdder neuron_2_add_1(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_1_p1), .Port2(neuron_2_add_1_p2), .Output_syn(neuron_2_add_1_out));
FixedPointAdder neuron_2_add_2(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_2_p1), .Port2(neuron_2_add_2_p2), .Output_syn(neuron_2_add_2_out));
FixedPointAdder neuron_2_add_3(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_3_p1), .Port2(neuron_2_add_3_p2), .Output_syn(neuron_2_add_3_out));
FixedPointAdder neuron_2_add_4(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_4_p1), .Port2(neuron_2_add_4_p2), .Output_syn(neuron_2_add_4_out));
FixedPointAdder neuron_2_add_5(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_5_p1), .Port2(neuron_2_add_5_p2), .Output_syn(neuron_2_add_5_out));
FixedPointAdder neuron_2_add_6(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_6_p1), .Port2(neuron_2_add_6_p2), .Output_syn(neuron_2_add_6_out));
FixedPointAdder neuron_2_add_7(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_7_p1), .Port2(neuron_2_add_7_p2), .Output_syn(neuron_2_add_7_out));
FixedPointAdder neuron_2_add_8(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_8_p1), .Port2(neuron_2_add_8_p2), .Output_syn(neuron_2_add_8_out));
FixedPointAdder neuron_2_add_9(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_9_p1), .Port2(neuron_2_add_9_p2), .Output_syn(neuron_2_add_9_out));
FixedPointAdder neuron_2_add_10(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_10_p1), .Port2(neuron_2_add_10_p2), .Output_syn(neuron_2_add_10_out));
FixedPointAdder neuron_2_add_11(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_11_p1), .Port2(neuron_2_add_11_p2), .Output_syn(neuron_2_add_11_out));
FixedPointAdder neuron_2_add_12(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_12_p1), .Port2(neuron_2_add_12_p2), .Output_syn(neuron_2_add_12_out));
FixedPointAdder neuron_2_add_13(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_13_p1), .Port2(neuron_2_add_13_p2), .Output_syn(neuron_2_add_13_out));
FixedPointAdder neuron_2_add_14(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_14_p1), .Port2(neuron_2_add_14_p2), .Output_syn(neuron_2_add_14_out));
FixedPointAdder neuron_2_add_15(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_15_p1), .Port2(neuron_2_add_15_p2), .Output_syn(neuron_2_add_15_out));
FixedPointAdder neuron_2_add_16(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_16_p1), .Port2(neuron_2_add_16_p2), .Output_syn(neuron_2_add_16_out));
FixedPointAdder neuron_2_add_17(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_17_p1), .Port2(neuron_2_add_17_p2), .Output_syn(neuron_2_add_17_out));
FixedPointAdder neuron_2_add_18(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_18_p1), .Port2(neuron_2_add_18_p2), .Output_syn(neuron_2_add_18_out));
FixedPointAdder neuron_2_add_19(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_19_p1), .Port2(neuron_2_add_19_p2), .Output_syn(neuron_2_add_19_out));
FixedPointAdder neuron_2_add_20(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_20_p1), .Port2(neuron_2_add_20_p2), .Output_syn(neuron_2_add_20_out));
FixedPointAdder neuron_2_add_21(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_21_p1), .Port2(neuron_2_add_21_p2), .Output_syn(neuron_2_add_21_out));
FixedPointAdder neuron_2_add_22(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_22_p1), .Port2(neuron_2_add_22_p2), .Output_syn(neuron_2_add_22_out));
FixedPointAdder neuron_2_add_23(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_23_p1), .Port2(neuron_2_add_23_p2), .Output_syn(neuron_2_add_23_out));
FixedPointAdder neuron_2_add_24(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_24_p1), .Port2(neuron_2_add_24_p2), .Output_syn(neuron_2_add_24_out));
FixedPointAdder neuron_2_add_25(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_25_p1), .Port2(neuron_2_add_25_p2), .Output_syn(neuron_2_add_25_out));
FixedPointAdder neuron_2_add_26(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_26_p1), .Port2(neuron_2_add_26_p2), .Output_syn(neuron_2_add_26_out));
FixedPointAdder neuron_2_add_27(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_2_add_27_p1), .Port2(neuron_2_add_27_p2), .Output_syn(neuron_2_add_27_out));

// neuron 3
FixedPointAdder neuron_3_add_0(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_0_p1), .Port2(neuron_3_add_0_p2), .Output_syn(neuron_3_add_0_out));
FixedPointAdder neuron_3_add_1(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_1_p1), .Port2(neuron_3_add_1_p2), .Output_syn(neuron_3_add_1_out));
FixedPointAdder neuron_3_add_2(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_2_p1), .Port2(neuron_3_add_2_p2), .Output_syn(neuron_3_add_2_out));
FixedPointAdder neuron_3_add_3(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_3_p1), .Port2(neuron_3_add_3_p2), .Output_syn(neuron_3_add_3_out));
FixedPointAdder neuron_3_add_4(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_4_p1), .Port2(neuron_3_add_4_p2), .Output_syn(neuron_3_add_4_out));
FixedPointAdder neuron_3_add_5(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_5_p1), .Port2(neuron_3_add_5_p2), .Output_syn(neuron_3_add_5_out));
FixedPointAdder neuron_3_add_6(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_6_p1), .Port2(neuron_3_add_6_p2), .Output_syn(neuron_3_add_6_out));
FixedPointAdder neuron_3_add_7(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_7_p1), .Port2(neuron_3_add_7_p2), .Output_syn(neuron_3_add_7_out));
FixedPointAdder neuron_3_add_8(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_8_p1), .Port2(neuron_3_add_8_p2), .Output_syn(neuron_3_add_8_out));
FixedPointAdder neuron_3_add_9(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_9_p1), .Port2(neuron_3_add_9_p2), .Output_syn(neuron_3_add_9_out));
FixedPointAdder neuron_3_add_10(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_10_p1), .Port2(neuron_3_add_10_p2), .Output_syn(neuron_3_add_10_out));
FixedPointAdder neuron_3_add_11(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_11_p1), .Port2(neuron_3_add_11_p2), .Output_syn(neuron_3_add_11_out));
FixedPointAdder neuron_3_add_12(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_12_p1), .Port2(neuron_3_add_12_p2), .Output_syn(neuron_3_add_12_out));
FixedPointAdder neuron_3_add_13(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_13_p1), .Port2(neuron_3_add_13_p2), .Output_syn(neuron_3_add_13_out));
FixedPointAdder neuron_3_add_14(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_14_p1), .Port2(neuron_3_add_14_p2), .Output_syn(neuron_3_add_14_out));
FixedPointAdder neuron_3_add_15(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_15_p1), .Port2(neuron_3_add_15_p2), .Output_syn(neuron_3_add_15_out));
FixedPointAdder neuron_3_add_16(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_16_p1), .Port2(neuron_3_add_16_p2), .Output_syn(neuron_3_add_16_out));
FixedPointAdder neuron_3_add_17(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_17_p1), .Port2(neuron_3_add_17_p2), .Output_syn(neuron_3_add_17_out));
FixedPointAdder neuron_3_add_18(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_18_p1), .Port2(neuron_3_add_18_p2), .Output_syn(neuron_3_add_18_out));
FixedPointAdder neuron_3_add_19(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_19_p1), .Port2(neuron_3_add_19_p2), .Output_syn(neuron_3_add_19_out));
FixedPointAdder neuron_3_add_20(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_20_p1), .Port2(neuron_3_add_20_p2), .Output_syn(neuron_3_add_20_out));
FixedPointAdder neuron_3_add_21(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_21_p1), .Port2(neuron_3_add_21_p2), .Output_syn(neuron_3_add_21_out));
FixedPointAdder neuron_3_add_22(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_22_p1), .Port2(neuron_3_add_22_p2), .Output_syn(neuron_3_add_22_out));
FixedPointAdder neuron_3_add_23(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_23_p1), .Port2(neuron_3_add_23_p2), .Output_syn(neuron_3_add_23_out));
FixedPointAdder neuron_3_add_24(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_24_p1), .Port2(neuron_3_add_24_p2), .Output_syn(neuron_3_add_24_out));
FixedPointAdder neuron_3_add_25(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_25_p1), .Port2(neuron_3_add_25_p2), .Output_syn(neuron_3_add_25_out));
FixedPointAdder neuron_3_add_26(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_26_p1), .Port2(neuron_3_add_26_p2), .Output_syn(neuron_3_add_26_out));
FixedPointAdder neuron_3_add_27(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_3_add_27_p1), .Port2(neuron_3_add_27_p2), .Output_syn(neuron_3_add_27_out));

// neuron 4
FixedPointAdder neuron_4_add_0(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_0_p1), .Port2(neuron_4_add_0_p2), .Output_syn(neuron_4_add_0_out));
FixedPointAdder neuron_4_add_1(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_1_p1), .Port2(neuron_4_add_1_p2), .Output_syn(neuron_4_add_1_out));
FixedPointAdder neuron_4_add_2(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_2_p1), .Port2(neuron_4_add_2_p2), .Output_syn(neuron_4_add_2_out));
FixedPointAdder neuron_4_add_3(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_3_p1), .Port2(neuron_4_add_3_p2), .Output_syn(neuron_4_add_3_out));
FixedPointAdder neuron_4_add_4(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_4_p1), .Port2(neuron_4_add_4_p2), .Output_syn(neuron_4_add_4_out));
FixedPointAdder neuron_4_add_5(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_5_p1), .Port2(neuron_4_add_5_p2), .Output_syn(neuron_4_add_5_out));
FixedPointAdder neuron_4_add_6(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_6_p1), .Port2(neuron_4_add_6_p2), .Output_syn(neuron_4_add_6_out));
FixedPointAdder neuron_4_add_7(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_7_p1), .Port2(neuron_4_add_7_p2), .Output_syn(neuron_4_add_7_out));
FixedPointAdder neuron_4_add_8(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_8_p1), .Port2(neuron_4_add_8_p2), .Output_syn(neuron_4_add_8_out));
FixedPointAdder neuron_4_add_9(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_9_p1), .Port2(neuron_4_add_9_p2), .Output_syn(neuron_4_add_9_out));
FixedPointAdder neuron_4_add_10(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_10_p1), .Port2(neuron_4_add_10_p2), .Output_syn(neuron_4_add_10_out));
FixedPointAdder neuron_4_add_11(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_11_p1), .Port2(neuron_4_add_11_p2), .Output_syn(neuron_4_add_11_out));
FixedPointAdder neuron_4_add_12(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_12_p1), .Port2(neuron_4_add_12_p2), .Output_syn(neuron_4_add_12_out));
FixedPointAdder neuron_4_add_13(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_13_p1), .Port2(neuron_4_add_13_p2), .Output_syn(neuron_4_add_13_out));
FixedPointAdder neuron_4_add_14(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_14_p1), .Port2(neuron_4_add_14_p2), .Output_syn(neuron_4_add_14_out));
FixedPointAdder neuron_4_add_15(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_15_p1), .Port2(neuron_4_add_15_p2), .Output_syn(neuron_4_add_15_out));
FixedPointAdder neuron_4_add_16(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_16_p1), .Port2(neuron_4_add_16_p2), .Output_syn(neuron_4_add_16_out));
FixedPointAdder neuron_4_add_17(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_17_p1), .Port2(neuron_4_add_17_p2), .Output_syn(neuron_4_add_17_out));
FixedPointAdder neuron_4_add_18(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_18_p1), .Port2(neuron_4_add_18_p2), .Output_syn(neuron_4_add_18_out));
FixedPointAdder neuron_4_add_19(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_19_p1), .Port2(neuron_4_add_19_p2), .Output_syn(neuron_4_add_19_out));
FixedPointAdder neuron_4_add_20(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_20_p1), .Port2(neuron_4_add_20_p2), .Output_syn(neuron_4_add_20_out));
FixedPointAdder neuron_4_add_21(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_21_p1), .Port2(neuron_4_add_21_p2), .Output_syn(neuron_4_add_21_out));
FixedPointAdder neuron_4_add_22(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_22_p1), .Port2(neuron_4_add_22_p2), .Output_syn(neuron_4_add_22_out));
FixedPointAdder neuron_4_add_23(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_23_p1), .Port2(neuron_4_add_23_p2), .Output_syn(neuron_4_add_23_out));
FixedPointAdder neuron_4_add_24(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_24_p1), .Port2(neuron_4_add_24_p2), .Output_syn(neuron_4_add_24_out));
FixedPointAdder neuron_4_add_25(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_25_p1), .Port2(neuron_4_add_25_p2), .Output_syn(neuron_4_add_25_out));
FixedPointAdder neuron_4_add_26(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_26_p1), .Port2(neuron_4_add_26_p2), .Output_syn(neuron_4_add_26_out));
FixedPointAdder neuron_4_add_27(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_4_add_27_p1), .Port2(neuron_4_add_27_p2), .Output_syn(neuron_4_add_27_out));

// neuron 5
FixedPointAdder neuron_5_add_0(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_0_p1), .Port2(neuron_5_add_0_p2), .Output_syn(neuron_5_add_0_out));
FixedPointAdder neuron_5_add_1(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_1_p1), .Port2(neuron_5_add_1_p2), .Output_syn(neuron_5_add_1_out));
FixedPointAdder neuron_5_add_2(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_2_p1), .Port2(neuron_5_add_2_p2), .Output_syn(neuron_5_add_2_out));
FixedPointAdder neuron_5_add_3(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_3_p1), .Port2(neuron_5_add_3_p2), .Output_syn(neuron_5_add_3_out));
FixedPointAdder neuron_5_add_4(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_4_p1), .Port2(neuron_5_add_4_p2), .Output_syn(neuron_5_add_4_out));
FixedPointAdder neuron_5_add_5(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_5_p1), .Port2(neuron_5_add_5_p2), .Output_syn(neuron_5_add_5_out));
FixedPointAdder neuron_5_add_6(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_6_p1), .Port2(neuron_5_add_6_p2), .Output_syn(neuron_5_add_6_out));
FixedPointAdder neuron_5_add_7(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_7_p1), .Port2(neuron_5_add_7_p2), .Output_syn(neuron_5_add_7_out));
FixedPointAdder neuron_5_add_8(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_8_p1), .Port2(neuron_5_add_8_p2), .Output_syn(neuron_5_add_8_out));
FixedPointAdder neuron_5_add_9(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_9_p1), .Port2(neuron_5_add_9_p2), .Output_syn(neuron_5_add_9_out));
FixedPointAdder neuron_5_add_10(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_10_p1), .Port2(neuron_5_add_10_p2), .Output_syn(neuron_5_add_10_out));
FixedPointAdder neuron_5_add_11(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_11_p1), .Port2(neuron_5_add_11_p2), .Output_syn(neuron_5_add_11_out));
FixedPointAdder neuron_5_add_12(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_12_p1), .Port2(neuron_5_add_12_p2), .Output_syn(neuron_5_add_12_out));
FixedPointAdder neuron_5_add_13(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_13_p1), .Port2(neuron_5_add_13_p2), .Output_syn(neuron_5_add_13_out));
FixedPointAdder neuron_5_add_14(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_14_p1), .Port2(neuron_5_add_14_p2), .Output_syn(neuron_5_add_14_out));
FixedPointAdder neuron_5_add_15(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_15_p1), .Port2(neuron_5_add_15_p2), .Output_syn(neuron_5_add_15_out));
FixedPointAdder neuron_5_add_16(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_16_p1), .Port2(neuron_5_add_16_p2), .Output_syn(neuron_5_add_16_out));
FixedPointAdder neuron_5_add_17(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_17_p1), .Port2(neuron_5_add_17_p2), .Output_syn(neuron_5_add_17_out));
FixedPointAdder neuron_5_add_18(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_18_p1), .Port2(neuron_5_add_18_p2), .Output_syn(neuron_5_add_18_out));
FixedPointAdder neuron_5_add_19(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_19_p1), .Port2(neuron_5_add_19_p2), .Output_syn(neuron_5_add_19_out));
FixedPointAdder neuron_5_add_20(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_20_p1), .Port2(neuron_5_add_20_p2), .Output_syn(neuron_5_add_20_out));
FixedPointAdder neuron_5_add_21(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_21_p1), .Port2(neuron_5_add_21_p2), .Output_syn(neuron_5_add_21_out));
FixedPointAdder neuron_5_add_22(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_22_p1), .Port2(neuron_5_add_22_p2), .Output_syn(neuron_5_add_22_out));
FixedPointAdder neuron_5_add_23(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_23_p1), .Port2(neuron_5_add_23_p2), .Output_syn(neuron_5_add_23_out));
FixedPointAdder neuron_5_add_24(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_24_p1), .Port2(neuron_5_add_24_p2), .Output_syn(neuron_5_add_24_out));
FixedPointAdder neuron_5_add_25(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_25_p1), .Port2(neuron_5_add_25_p2), .Output_syn(neuron_5_add_25_out));
FixedPointAdder neuron_5_add_26(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_26_p1), .Port2(neuron_5_add_26_p2), .Output_syn(neuron_5_add_26_out));
FixedPointAdder neuron_5_add_27(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_5_add_27_p1), .Port2(neuron_5_add_27_p2), .Output_syn(neuron_5_add_27_out));

// neuron 6
FixedPointAdder neuron_6_add_0(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_0_p1), .Port2(neuron_6_add_0_p2), .Output_syn(neuron_6_add_0_out));
FixedPointAdder neuron_6_add_1(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_1_p1), .Port2(neuron_6_add_1_p2), .Output_syn(neuron_6_add_1_out));
FixedPointAdder neuron_6_add_2(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_2_p1), .Port2(neuron_6_add_2_p2), .Output_syn(neuron_6_add_2_out));
FixedPointAdder neuron_6_add_3(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_3_p1), .Port2(neuron_6_add_3_p2), .Output_syn(neuron_6_add_3_out));
FixedPointAdder neuron_6_add_4(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_4_p1), .Port2(neuron_6_add_4_p2), .Output_syn(neuron_6_add_4_out));
FixedPointAdder neuron_6_add_5(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_5_p1), .Port2(neuron_6_add_5_p2), .Output_syn(neuron_6_add_5_out));
FixedPointAdder neuron_6_add_6(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_6_p1), .Port2(neuron_6_add_6_p2), .Output_syn(neuron_6_add_6_out));
FixedPointAdder neuron_6_add_7(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_7_p1), .Port2(neuron_6_add_7_p2), .Output_syn(neuron_6_add_7_out));
FixedPointAdder neuron_6_add_8(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_8_p1), .Port2(neuron_6_add_8_p2), .Output_syn(neuron_6_add_8_out));
FixedPointAdder neuron_6_add_9(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_9_p1), .Port2(neuron_6_add_9_p2), .Output_syn(neuron_6_add_9_out));
FixedPointAdder neuron_6_add_10(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_10_p1), .Port2(neuron_6_add_10_p2), .Output_syn(neuron_6_add_10_out));
FixedPointAdder neuron_6_add_11(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_11_p1), .Port2(neuron_6_add_11_p2), .Output_syn(neuron_6_add_11_out));
FixedPointAdder neuron_6_add_12(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_12_p1), .Port2(neuron_6_add_12_p2), .Output_syn(neuron_6_add_12_out));
FixedPointAdder neuron_6_add_13(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_13_p1), .Port2(neuron_6_add_13_p2), .Output_syn(neuron_6_add_13_out));
FixedPointAdder neuron_6_add_14(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_14_p1), .Port2(neuron_6_add_14_p2), .Output_syn(neuron_6_add_14_out));
FixedPointAdder neuron_6_add_15(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_15_p1), .Port2(neuron_6_add_15_p2), .Output_syn(neuron_6_add_15_out));
FixedPointAdder neuron_6_add_16(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_16_p1), .Port2(neuron_6_add_16_p2), .Output_syn(neuron_6_add_16_out));
FixedPointAdder neuron_6_add_17(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_17_p1), .Port2(neuron_6_add_17_p2), .Output_syn(neuron_6_add_17_out));
FixedPointAdder neuron_6_add_18(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_18_p1), .Port2(neuron_6_add_18_p2), .Output_syn(neuron_6_add_18_out));
FixedPointAdder neuron_6_add_19(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_19_p1), .Port2(neuron_6_add_19_p2), .Output_syn(neuron_6_add_19_out));
FixedPointAdder neuron_6_add_20(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_20_p1), .Port2(neuron_6_add_20_p2), .Output_syn(neuron_6_add_20_out));
FixedPointAdder neuron_6_add_21(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_21_p1), .Port2(neuron_6_add_21_p2), .Output_syn(neuron_6_add_21_out));
FixedPointAdder neuron_6_add_22(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_22_p1), .Port2(neuron_6_add_22_p2), .Output_syn(neuron_6_add_22_out));
FixedPointAdder neuron_6_add_23(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_23_p1), .Port2(neuron_6_add_23_p2), .Output_syn(neuron_6_add_23_out));
FixedPointAdder neuron_6_add_24(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_24_p1), .Port2(neuron_6_add_24_p2), .Output_syn(neuron_6_add_24_out));
FixedPointAdder neuron_6_add_25(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_25_p1), .Port2(neuron_6_add_25_p2), .Output_syn(neuron_6_add_25_out));
FixedPointAdder neuron_6_add_26(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_26_p1), .Port2(neuron_6_add_26_p2), .Output_syn(neuron_6_add_26_out));
FixedPointAdder neuron_6_add_27(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_6_add_27_p1), .Port2(neuron_6_add_27_p2), .Output_syn(neuron_6_add_27_out));

// neuron 7
FixedPointAdder neuron_7_add_0(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_0_p1), .Port2(neuron_7_add_0_p2), .Output_syn(neuron_7_add_0_out));
FixedPointAdder neuron_7_add_1(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_1_p1), .Port2(neuron_7_add_1_p2), .Output_syn(neuron_7_add_1_out));
FixedPointAdder neuron_7_add_2(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_2_p1), .Port2(neuron_7_add_2_p2), .Output_syn(neuron_7_add_2_out));
FixedPointAdder neuron_7_add_3(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_3_p1), .Port2(neuron_7_add_3_p2), .Output_syn(neuron_7_add_3_out));
FixedPointAdder neuron_7_add_4(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_4_p1), .Port2(neuron_7_add_4_p2), .Output_syn(neuron_7_add_4_out));
FixedPointAdder neuron_7_add_5(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_5_p1), .Port2(neuron_7_add_5_p2), .Output_syn(neuron_7_add_5_out));
FixedPointAdder neuron_7_add_6(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_6_p1), .Port2(neuron_7_add_6_p2), .Output_syn(neuron_7_add_6_out));
FixedPointAdder neuron_7_add_7(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_7_p1), .Port2(neuron_7_add_7_p2), .Output_syn(neuron_7_add_7_out));
FixedPointAdder neuron_7_add_8(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_8_p1), .Port2(neuron_7_add_8_p2), .Output_syn(neuron_7_add_8_out));
FixedPointAdder neuron_7_add_9(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_9_p1), .Port2(neuron_7_add_9_p2), .Output_syn(neuron_7_add_9_out));
FixedPointAdder neuron_7_add_10(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_10_p1), .Port2(neuron_7_add_10_p2), .Output_syn(neuron_7_add_10_out));
FixedPointAdder neuron_7_add_11(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_11_p1), .Port2(neuron_7_add_11_p2), .Output_syn(neuron_7_add_11_out));
FixedPointAdder neuron_7_add_12(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_12_p1), .Port2(neuron_7_add_12_p2), .Output_syn(neuron_7_add_12_out));
FixedPointAdder neuron_7_add_13(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_13_p1), .Port2(neuron_7_add_13_p2), .Output_syn(neuron_7_add_13_out));
FixedPointAdder neuron_7_add_14(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_14_p1), .Port2(neuron_7_add_14_p2), .Output_syn(neuron_7_add_14_out));
FixedPointAdder neuron_7_add_15(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_15_p1), .Port2(neuron_7_add_15_p2), .Output_syn(neuron_7_add_15_out));
FixedPointAdder neuron_7_add_16(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_16_p1), .Port2(neuron_7_add_16_p2), .Output_syn(neuron_7_add_16_out));
FixedPointAdder neuron_7_add_17(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_17_p1), .Port2(neuron_7_add_17_p2), .Output_syn(neuron_7_add_17_out));
FixedPointAdder neuron_7_add_18(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_18_p1), .Port2(neuron_7_add_18_p2), .Output_syn(neuron_7_add_18_out));
FixedPointAdder neuron_7_add_19(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_19_p1), .Port2(neuron_7_add_19_p2), .Output_syn(neuron_7_add_19_out));
FixedPointAdder neuron_7_add_20(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_20_p1), .Port2(neuron_7_add_20_p2), .Output_syn(neuron_7_add_20_out));
FixedPointAdder neuron_7_add_21(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_21_p1), .Port2(neuron_7_add_21_p2), .Output_syn(neuron_7_add_21_out));
FixedPointAdder neuron_7_add_22(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_22_p1), .Port2(neuron_7_add_22_p2), .Output_syn(neuron_7_add_22_out));
FixedPointAdder neuron_7_add_23(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_23_p1), .Port2(neuron_7_add_23_p2), .Output_syn(neuron_7_add_23_out));
FixedPointAdder neuron_7_add_24(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_24_p1), .Port2(neuron_7_add_24_p2), .Output_syn(neuron_7_add_24_out));
FixedPointAdder neuron_7_add_25(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_25_p1), .Port2(neuron_7_add_25_p2), .Output_syn(neuron_7_add_25_out));
FixedPointAdder neuron_7_add_26(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_26_p1), .Port2(neuron_7_add_26_p2), .Output_syn(neuron_7_add_26_out));
FixedPointAdder neuron_7_add_27(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_7_add_27_p1), .Port2(neuron_7_add_27_p2), .Output_syn(neuron_7_add_27_out));

// neuron 8
FixedPointAdder neuron_8_add_0(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_0_p1), .Port2(neuron_8_add_0_p2), .Output_syn(neuron_8_add_0_out));
FixedPointAdder neuron_8_add_1(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_1_p1), .Port2(neuron_8_add_1_p2), .Output_syn(neuron_8_add_1_out));
FixedPointAdder neuron_8_add_2(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_2_p1), .Port2(neuron_8_add_2_p2), .Output_syn(neuron_8_add_2_out));
FixedPointAdder neuron_8_add_3(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_3_p1), .Port2(neuron_8_add_3_p2), .Output_syn(neuron_8_add_3_out));
FixedPointAdder neuron_8_add_4(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_4_p1), .Port2(neuron_8_add_4_p2), .Output_syn(neuron_8_add_4_out));
FixedPointAdder neuron_8_add_5(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_5_p1), .Port2(neuron_8_add_5_p2), .Output_syn(neuron_8_add_5_out));
FixedPointAdder neuron_8_add_6(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_6_p1), .Port2(neuron_8_add_6_p2), .Output_syn(neuron_8_add_6_out));
FixedPointAdder neuron_8_add_7(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_7_p1), .Port2(neuron_8_add_7_p2), .Output_syn(neuron_8_add_7_out));
FixedPointAdder neuron_8_add_8(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_8_p1), .Port2(neuron_8_add_8_p2), .Output_syn(neuron_8_add_8_out));
FixedPointAdder neuron_8_add_9(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_9_p1), .Port2(neuron_8_add_9_p2), .Output_syn(neuron_8_add_9_out));
FixedPointAdder neuron_8_add_10(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_10_p1), .Port2(neuron_8_add_10_p2), .Output_syn(neuron_8_add_10_out));
FixedPointAdder neuron_8_add_11(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_11_p1), .Port2(neuron_8_add_11_p2), .Output_syn(neuron_8_add_11_out));
FixedPointAdder neuron_8_add_12(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_12_p1), .Port2(neuron_8_add_12_p2), .Output_syn(neuron_8_add_12_out));
FixedPointAdder neuron_8_add_13(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_13_p1), .Port2(neuron_8_add_13_p2), .Output_syn(neuron_8_add_13_out));
FixedPointAdder neuron_8_add_14(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_14_p1), .Port2(neuron_8_add_14_p2), .Output_syn(neuron_8_add_14_out));
FixedPointAdder neuron_8_add_15(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_15_p1), .Port2(neuron_8_add_15_p2), .Output_syn(neuron_8_add_15_out));
FixedPointAdder neuron_8_add_16(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_16_p1), .Port2(neuron_8_add_16_p2), .Output_syn(neuron_8_add_16_out));
FixedPointAdder neuron_8_add_17(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_17_p1), .Port2(neuron_8_add_17_p2), .Output_syn(neuron_8_add_17_out));
FixedPointAdder neuron_8_add_18(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_18_p1), .Port2(neuron_8_add_18_p2), .Output_syn(neuron_8_add_18_out));
FixedPointAdder neuron_8_add_19(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_19_p1), .Port2(neuron_8_add_19_p2), .Output_syn(neuron_8_add_19_out));
FixedPointAdder neuron_8_add_20(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_20_p1), .Port2(neuron_8_add_20_p2), .Output_syn(neuron_8_add_20_out));
FixedPointAdder neuron_8_add_21(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_21_p1), .Port2(neuron_8_add_21_p2), .Output_syn(neuron_8_add_21_out));
FixedPointAdder neuron_8_add_22(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_22_p1), .Port2(neuron_8_add_22_p2), .Output_syn(neuron_8_add_22_out));
FixedPointAdder neuron_8_add_23(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_23_p1), .Port2(neuron_8_add_23_p2), .Output_syn(neuron_8_add_23_out));
FixedPointAdder neuron_8_add_24(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_24_p1), .Port2(neuron_8_add_24_p2), .Output_syn(neuron_8_add_24_out));
FixedPointAdder neuron_8_add_25(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_25_p1), .Port2(neuron_8_add_25_p2), .Output_syn(neuron_8_add_25_out));
FixedPointAdder neuron_8_add_26(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_26_p1), .Port2(neuron_8_add_26_p2), .Output_syn(neuron_8_add_26_out));
FixedPointAdder neuron_8_add_27(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_8_add_27_p1), .Port2(neuron_8_add_27_p2), .Output_syn(neuron_8_add_27_out));

// neuron 9
FixedPointAdder neuron_9_add_0(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_0_p1), .Port2(neuron_9_add_0_p2), .Output_syn(neuron_9_add_0_out));
FixedPointAdder neuron_9_add_1(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_1_p1), .Port2(neuron_9_add_1_p2), .Output_syn(neuron_9_add_1_out));
FixedPointAdder neuron_9_add_2(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_2_p1), .Port2(neuron_9_add_2_p2), .Output_syn(neuron_9_add_2_out));
FixedPointAdder neuron_9_add_3(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_3_p1), .Port2(neuron_9_add_3_p2), .Output_syn(neuron_9_add_3_out));
FixedPointAdder neuron_9_add_4(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_4_p1), .Port2(neuron_9_add_4_p2), .Output_syn(neuron_9_add_4_out));
FixedPointAdder neuron_9_add_5(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_5_p1), .Port2(neuron_9_add_5_p2), .Output_syn(neuron_9_add_5_out));
FixedPointAdder neuron_9_add_6(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_6_p1), .Port2(neuron_9_add_6_p2), .Output_syn(neuron_9_add_6_out));
FixedPointAdder neuron_9_add_7(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_7_p1), .Port2(neuron_9_add_7_p2), .Output_syn(neuron_9_add_7_out));
FixedPointAdder neuron_9_add_8(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_8_p1), .Port2(neuron_9_add_8_p2), .Output_syn(neuron_9_add_8_out));
FixedPointAdder neuron_9_add_9(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_9_p1), .Port2(neuron_9_add_9_p2), .Output_syn(neuron_9_add_9_out));
FixedPointAdder neuron_9_add_10(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_10_p1), .Port2(neuron_9_add_10_p2), .Output_syn(neuron_9_add_10_out));
FixedPointAdder neuron_9_add_11(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_11_p1), .Port2(neuron_9_add_11_p2), .Output_syn(neuron_9_add_11_out));
FixedPointAdder neuron_9_add_12(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_12_p1), .Port2(neuron_9_add_12_p2), .Output_syn(neuron_9_add_12_out));
FixedPointAdder neuron_9_add_13(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_13_p1), .Port2(neuron_9_add_13_p2), .Output_syn(neuron_9_add_13_out));
FixedPointAdder neuron_9_add_14(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_14_p1), .Port2(neuron_9_add_14_p2), .Output_syn(neuron_9_add_14_out));
FixedPointAdder neuron_9_add_15(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_15_p1), .Port2(neuron_9_add_15_p2), .Output_syn(neuron_9_add_15_out));
FixedPointAdder neuron_9_add_16(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_16_p1), .Port2(neuron_9_add_16_p2), .Output_syn(neuron_9_add_16_out));
FixedPointAdder neuron_9_add_17(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_17_p1), .Port2(neuron_9_add_17_p2), .Output_syn(neuron_9_add_17_out));
FixedPointAdder neuron_9_add_18(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_18_p1), .Port2(neuron_9_add_18_p2), .Output_syn(neuron_9_add_18_out));
FixedPointAdder neuron_9_add_19(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_19_p1), .Port2(neuron_9_add_19_p2), .Output_syn(neuron_9_add_19_out));
FixedPointAdder neuron_9_add_20(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_20_p1), .Port2(neuron_9_add_20_p2), .Output_syn(neuron_9_add_20_out));
FixedPointAdder neuron_9_add_21(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_21_p1), .Port2(neuron_9_add_21_p2), .Output_syn(neuron_9_add_21_out));
FixedPointAdder neuron_9_add_22(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_22_p1), .Port2(neuron_9_add_22_p2), .Output_syn(neuron_9_add_22_out));
FixedPointAdder neuron_9_add_23(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_23_p1), .Port2(neuron_9_add_23_p2), .Output_syn(neuron_9_add_23_out));
FixedPointAdder neuron_9_add_24(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_24_p1), .Port2(neuron_9_add_24_p2), .Output_syn(neuron_9_add_24_out));
FixedPointAdder neuron_9_add_25(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_25_p1), .Port2(neuron_9_add_25_p2), .Output_syn(neuron_9_add_25_out));
FixedPointAdder neuron_9_add_26(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_26_p1), .Port2(neuron_9_add_26_p2), .Output_syn(neuron_9_add_26_out));
FixedPointAdder neuron_9_add_27(.clk(neuron_clk), .GlobalReset(globalreset), .Port1(neuron_9_add_27_p1), .Port2(neuron_9_add_27_p2), .Output_syn(neuron_9_add_27_out));

// Initialize input for neuron multiplier pixels
// Timing might need to be adjusted
Neuron_mul_pixel neuron_mul_pixel(
.neuron_clk,
.globalreset,
.N,
.Pix_0,.Pix_1,.Pix_2,.Pix_3,.Pix_4,.Pix_5,.Pix_6,.Pix_7,.Pix_8,.Pix_9,.Pix_10,.Pix_11,.Pix_12,.Pix_13,.Pix_14,.Pix_15,.Pix_16,.Pix_17,.Pix_18,.Pix_19,.Pix_20,.Pix_21,.Pix_22,.Pix_23,.Pix_24,.Pix_25,.Pix_26,.Pix_27,.Pix_28,.Pix_29,.Pix_30,.Pix_31,.Pix_32,.Pix_33,.Pix_34,.Pix_35,.Pix_36,.Pix_37,.Pix_38,.Pix_39,.Pix_40,.Pix_41,.Pix_42,.Pix_43,.Pix_44,.Pix_45,.Pix_46,.Pix_47,.Pix_48,.Pix_49,.Pix_50,.Pix_51,.Pix_52,.Pix_53,.Pix_54,.Pix_55,.Pix_56,.Pix_57,.Pix_58,.Pix_59,.Pix_60,.Pix_61,.Pix_62,.Pix_63,.Pix_64,.Pix_65,.Pix_66,.Pix_67,.Pix_68,.Pix_69,.Pix_70,.Pix_71,.Pix_72,.Pix_73,.Pix_74,.Pix_75,.Pix_76,.Pix_77,.Pix_78,.Pix_79,.Pix_80,.Pix_81,.Pix_82,.Pix_83,.Pix_84,.Pix_85,.Pix_86,.Pix_87,.Pix_88,.Pix_89,.Pix_90,.Pix_91,.Pix_92,.Pix_93,.Pix_94,.Pix_95,.Pix_96,.Pix_97,.Pix_98,.Pix_99,.Pix_100,.Pix_101,.Pix_102,.Pix_103,.Pix_104,.Pix_105,.Pix_106,.Pix_107,.Pix_108,.Pix_109,.Pix_110,.Pix_111,.Pix_112,.Pix_113,.Pix_114,.Pix_115,.Pix_116,.Pix_117,.Pix_118,.Pix_119,.Pix_120,.Pix_121,.Pix_122,.Pix_123,.Pix_124,.Pix_125,.Pix_126,.Pix_127,.Pix_128,.Pix_129,.Pix_130,.Pix_131,.Pix_132,.Pix_133,.Pix_134,.Pix_135,.Pix_136,.Pix_137,.Pix_138,.Pix_139,.Pix_140,.Pix_141,.Pix_142,.Pix_143,.Pix_144,.Pix_145,.Pix_146,.Pix_147,.Pix_148,.Pix_149,.Pix_150,.Pix_151,.Pix_152,.Pix_153,.Pix_154,.Pix_155,.Pix_156,.Pix_157,.Pix_158,.Pix_159,.Pix_160,.Pix_161,.Pix_162,.Pix_163,.Pix_164,.Pix_165,.Pix_166,.Pix_167,.Pix_168,.Pix_169,.Pix_170,.Pix_171,.Pix_172,.Pix_173,.Pix_174,.Pix_175,.Pix_176,.Pix_177,.Pix_178,.Pix_179,.Pix_180,.Pix_181,.Pix_182,.Pix_183,.Pix_184,.Pix_185,.Pix_186,.Pix_187,.Pix_188,.Pix_189,.Pix_190,.Pix_191,.Pix_192,.Pix_193,.Pix_194,.Pix_195,.Pix_196,.Pix_197,.Pix_198,.Pix_199,.Pix_200,.Pix_201,.Pix_202,.Pix_203,.Pix_204,.Pix_205,.Pix_206,.Pix_207,.Pix_208,.Pix_209,.Pix_210,.Pix_211,.Pix_212,.Pix_213,.Pix_214,.Pix_215,.Pix_216,.Pix_217,.Pix_218,.Pix_219,.Pix_220,.Pix_221,.Pix_222,.Pix_223,.Pix_224,.Pix_225,.Pix_226,.Pix_227,.Pix_228,.Pix_229,.Pix_230,.Pix_231,.Pix_232,.Pix_233,.Pix_234,.Pix_235,.Pix_236,.Pix_237,.Pix_238,.Pix_239,.Pix_240,.Pix_241,.Pix_242,.Pix_243,.Pix_244,.Pix_245,.Pix_246,.Pix_247,.Pix_248,.Pix_249,.Pix_250,.Pix_251,.Pix_252,.Pix_253,.Pix_254,.Pix_255,.Pix_256,.Pix_257,.Pix_258,.Pix_259,.Pix_260,.Pix_261,.Pix_262,.Pix_263,.Pix_264,.Pix_265,.Pix_266,.Pix_267,.Pix_268,.Pix_269,.Pix_270,.Pix_271,.Pix_272,.Pix_273,.Pix_274,.Pix_275,.Pix_276,.Pix_277,.Pix_278,.Pix_279,.Pix_280,.Pix_281,.Pix_282,.Pix_283,.Pix_284,.Pix_285,.Pix_286,.Pix_287,.Pix_288,.Pix_289,.Pix_290,.Pix_291,.Pix_292,.Pix_293,.Pix_294,.Pix_295,.Pix_296,.Pix_297,.Pix_298,.Pix_299,.Pix_300,.Pix_301,.Pix_302,.Pix_303,.Pix_304,.Pix_305,.Pix_306,.Pix_307,.Pix_308,.Pix_309,.Pix_310,.Pix_311,.Pix_312,.Pix_313,.Pix_314,.Pix_315,.Pix_316,.Pix_317,.Pix_318,.Pix_319,.Pix_320,.Pix_321,.Pix_322,.Pix_323,.Pix_324,.Pix_325,.Pix_326,.Pix_327,.Pix_328,.Pix_329,.Pix_330,.Pix_331,.Pix_332,.Pix_333,.Pix_334,.Pix_335,.Pix_336,.Pix_337,.Pix_338,.Pix_339,.Pix_340,.Pix_341,.Pix_342,.Pix_343,.Pix_344,.Pix_345,.Pix_346,.Pix_347,.Pix_348,.Pix_349,.Pix_350,.Pix_351,.Pix_352,.Pix_353,.Pix_354,.Pix_355,.Pix_356,.Pix_357,.Pix_358,.Pix_359,.Pix_360,.Pix_361,.Pix_362,.Pix_363,.Pix_364,.Pix_365,.Pix_366,.Pix_367,.Pix_368,.Pix_369,.Pix_370,.Pix_371,.Pix_372,.Pix_373,.Pix_374,.Pix_375,.Pix_376,.Pix_377,.Pix_378,.Pix_379,.Pix_380,.Pix_381,.Pix_382,.Pix_383,.Pix_384,.Pix_385,.Pix_386,.Pix_387,.Pix_388,.Pix_389,.Pix_390,.Pix_391,.Pix_392,.Pix_393,.Pix_394,.Pix_395,.Pix_396,.Pix_397,.Pix_398,.Pix_399,.Pix_400,.Pix_401,.Pix_402,.Pix_403,.Pix_404,.Pix_405,.Pix_406,.Pix_407,.Pix_408,.Pix_409,.Pix_410,.Pix_411,.Pix_412,.Pix_413,.Pix_414,.Pix_415,.Pix_416,.Pix_417,.Pix_418,.Pix_419,.Pix_420,.Pix_421,.Pix_422,.Pix_423,.Pix_424,.Pix_425,.Pix_426,.Pix_427,.Pix_428,.Pix_429,.Pix_430,.Pix_431,.Pix_432,.Pix_433,.Pix_434,.Pix_435,.Pix_436,.Pix_437,.Pix_438,.Pix_439,.Pix_440,.Pix_441,.Pix_442,.Pix_443,.Pix_444,.Pix_445,.Pix_446,.Pix_447,.Pix_448,.Pix_449,.Pix_450,.Pix_451,.Pix_452,.Pix_453,.Pix_454,.Pix_455,.Pix_456,.Pix_457,.Pix_458,.Pix_459,.Pix_460,.Pix_461,.Pix_462,.Pix_463,.Pix_464,.Pix_465,.Pix_466,.Pix_467,.Pix_468,.Pix_469,.Pix_470,.Pix_471,.Pix_472,.Pix_473,.Pix_474,.Pix_475,.Pix_476,.Pix_477,.Pix_478,.Pix_479,.Pix_480,.Pix_481,.Pix_482,.Pix_483,.Pix_484,.Pix_485,.Pix_486,.Pix_487,.Pix_488,.Pix_489,.Pix_490,.Pix_491,.Pix_492,.Pix_493,.Pix_494,.Pix_495,.Pix_496,.Pix_497,.Pix_498,.Pix_499,.Pix_500,.Pix_501,.Pix_502,.Pix_503,.Pix_504,.Pix_505,.Pix_506,.Pix_507,.Pix_508,.Pix_509,.Pix_510,.Pix_511,.Pix_512,.Pix_513,.Pix_514,.Pix_515,.Pix_516,.Pix_517,.Pix_518,.Pix_519,.Pix_520,.Pix_521,.Pix_522,.Pix_523,.Pix_524,.Pix_525,.Pix_526,.Pix_527,.Pix_528,.Pix_529,.Pix_530,.Pix_531,.Pix_532,.Pix_533,.Pix_534,.Pix_535,.Pix_536,.Pix_537,.Pix_538,.Pix_539,.Pix_540,.Pix_541,.Pix_542,.Pix_543,.Pix_544,.Pix_545,.Pix_546,.Pix_547,.Pix_548,.Pix_549,.Pix_550,.Pix_551,.Pix_552,.Pix_553,.Pix_554,.Pix_555,.Pix_556,.Pix_557,.Pix_558,.Pix_559,.Pix_560,.Pix_561,.Pix_562,.Pix_563,.Pix_564,.Pix_565,.Pix_566,.Pix_567,.Pix_568,.Pix_569,.Pix_570,.Pix_571,.Pix_572,.Pix_573,.Pix_574,.Pix_575,.Pix_576,.Pix_577,.Pix_578,.Pix_579,.Pix_580,.Pix_581,.Pix_582,.Pix_583,.Pix_584,.Pix_585,.Pix_586,.Pix_587,.Pix_588,.Pix_589,.Pix_590,.Pix_591,.Pix_592,.Pix_593,.Pix_594,.Pix_595,.Pix_596,.Pix_597,.Pix_598,.Pix_599,.Pix_600,.Pix_601,.Pix_602,.Pix_603,.Pix_604,.Pix_605,.Pix_606,.Pix_607,.Pix_608,.Pix_609,.Pix_610,.Pix_611,.Pix_612,.Pix_613,.Pix_614,.Pix_615,.Pix_616,.Pix_617,.Pix_618,.Pix_619,.Pix_620,.Pix_621,.Pix_622,.Pix_623,.Pix_624,.Pix_625,.Pix_626,.Pix_627,.Pix_628,.Pix_629,.Pix_630,.Pix_631,.Pix_632,.Pix_633,.Pix_634,.Pix_635,.Pix_636,.Pix_637,.Pix_638,.Pix_639,.Pix_640,.Pix_641,.Pix_642,.Pix_643,.Pix_644,.Pix_645,.Pix_646,.Pix_647,.Pix_648,.Pix_649,.Pix_650,.Pix_651,.Pix_652,.Pix_653,.Pix_654,.Pix_655,.Pix_656,.Pix_657,.Pix_658,.Pix_659,.Pix_660,.Pix_661,.Pix_662,.Pix_663,.Pix_664,.Pix_665,.Pix_666,.Pix_667,.Pix_668,.Pix_669,.Pix_670,.Pix_671,.Pix_672,.Pix_673,.Pix_674,.Pix_675,.Pix_676,.Pix_677,.Pix_678,.Pix_679,.Pix_680,.Pix_681,.Pix_682,.Pix_683,.Pix_684,.Pix_685,.Pix_686,.Pix_687,.Pix_688,.Pix_689,.Pix_690,.Pix_691,.Pix_692,.Pix_693,.Pix_694,.Pix_695,.Pix_696,.Pix_697,.Pix_698,.Pix_699,.Pix_700,.Pix_701,.Pix_702,.Pix_703,.Pix_704,.Pix_705,.Pix_706,.Pix_707,.Pix_708,.Pix_709,.Pix_710,.Pix_711,.Pix_712,.Pix_713,.Pix_714,.Pix_715,.Pix_716,.Pix_717,.Pix_718,.Pix_719,.Pix_720,.Pix_721,.Pix_722,.Pix_723,.Pix_724,.Pix_725,.Pix_726,.Pix_727,.Pix_728,.Pix_729,.Pix_730,.Pix_731,.Pix_732,.Pix_733,.Pix_734,.Pix_735,.Pix_736,.Pix_737,.Pix_738,.Pix_739,.Pix_740,.Pix_741,.Pix_742,.Pix_743,.Pix_744,.Pix_745,.Pix_746,.Pix_747,.Pix_748,.Pix_749,.Pix_750,.Pix_751,.Pix_752,.Pix_753,.Pix_754,.Pix_755,.Pix_756,.Pix_757,.Pix_758,.Pix_759,.Pix_760,.Pix_761,.Pix_762,.Pix_763,.Pix_764,.Pix_765,.Pix_766,.Pix_767,.Pix_768,.Pix_769,.Pix_770,.Pix_771,.Pix_772,.Pix_773,.Pix_774,.Pix_775,.Pix_776,.Pix_777,.Pix_778,.Pix_779,.Pix_780,.Pix_781,.Pix_782,.Pix_783,.Pix_784,
.neuron_mul_0_p, .neuron_mul_1_p, .neuron_mul_2_p, .neuron_mul_3_p, .neuron_mul_4_p, .neuron_mul_5_p, .neuron_mul_6_p, .neuron_mul_7_p, .neuron_mul_8_p, .neuron_mul_9_p, .neuron_mul_10_p, .neuron_mul_11_p, .neuron_mul_12_p, .neuron_mul_13_p, .neuron_mul_14_p, .neuron_mul_15_p, .neuron_mul_16_p, .neuron_mul_17_p, .neuron_mul_18_p, .neuron_mul_19_p, .neuron_mul_20_p, .neuron_mul_21_p, .neuron_mul_22_p, .neuron_mul_23_p, .neuron_mul_24_p, .neuron_mul_25_p, .neuron_mul_26_p, .neuron_mul_27_p
);

Neuron_mul_weight neuron_mul_weight(
.neuron_clk,
.globalreset,
.N,
.Wgt_0_0,.Wgt_0_1,.Wgt_0_2,.Wgt_0_3,.Wgt_0_4,.Wgt_0_5,.Wgt_0_6,.Wgt_0_7,.Wgt_0_8,.Wgt_0_9,.Wgt_0_10,.Wgt_0_11,.Wgt_0_12,.Wgt_0_13,.Wgt_0_14,.Wgt_0_15,.Wgt_0_16,.Wgt_0_17,.Wgt_0_18,.Wgt_0_19,.Wgt_0_20,.Wgt_0_21,.Wgt_0_22,.Wgt_0_23,.Wgt_0_24,.Wgt_0_25,.Wgt_0_26,.Wgt_0_27,.Wgt_0_28,.Wgt_0_29,.Wgt_0_30,.Wgt_0_31,.Wgt_0_32,.Wgt_0_33,.Wgt_0_34,.Wgt_0_35,.Wgt_0_36,.Wgt_0_37,.Wgt_0_38,.Wgt_0_39,.Wgt_0_40,.Wgt_0_41,.Wgt_0_42,.Wgt_0_43,.Wgt_0_44,.Wgt_0_45,.Wgt_0_46,.Wgt_0_47,.Wgt_0_48,.Wgt_0_49,.Wgt_0_50,.Wgt_0_51,.Wgt_0_52,.Wgt_0_53,.Wgt_0_54,.Wgt_0_55,.Wgt_0_56,.Wgt_0_57,.Wgt_0_58,.Wgt_0_59,.Wgt_0_60,.Wgt_0_61,.Wgt_0_62,.Wgt_0_63,.Wgt_0_64,.Wgt_0_65,.Wgt_0_66,.Wgt_0_67,.Wgt_0_68,.Wgt_0_69,.Wgt_0_70,.Wgt_0_71,.Wgt_0_72,.Wgt_0_73,.Wgt_0_74,.Wgt_0_75,.Wgt_0_76,.Wgt_0_77,.Wgt_0_78,.Wgt_0_79,.Wgt_0_80,.Wgt_0_81,.Wgt_0_82,.Wgt_0_83,.Wgt_0_84,.Wgt_0_85,.Wgt_0_86,.Wgt_0_87,.Wgt_0_88,.Wgt_0_89,.Wgt_0_90,.Wgt_0_91,.Wgt_0_92,.Wgt_0_93,.Wgt_0_94,.Wgt_0_95,.Wgt_0_96,.Wgt_0_97,.Wgt_0_98,.Wgt_0_99,.Wgt_0_100,.Wgt_0_101,.Wgt_0_102,.Wgt_0_103,.Wgt_0_104,.Wgt_0_105,.Wgt_0_106,.Wgt_0_107,.Wgt_0_108,.Wgt_0_109,.Wgt_0_110,.Wgt_0_111,.Wgt_0_112,.Wgt_0_113,.Wgt_0_114,.Wgt_0_115,.Wgt_0_116,.Wgt_0_117,.Wgt_0_118,.Wgt_0_119,.Wgt_0_120,.Wgt_0_121,.Wgt_0_122,.Wgt_0_123,.Wgt_0_124,.Wgt_0_125,.Wgt_0_126,.Wgt_0_127,.Wgt_0_128,.Wgt_0_129,.Wgt_0_130,.Wgt_0_131,.Wgt_0_132,.Wgt_0_133,.Wgt_0_134,.Wgt_0_135,.Wgt_0_136,.Wgt_0_137,.Wgt_0_138,.Wgt_0_139,.Wgt_0_140,.Wgt_0_141,.Wgt_0_142,.Wgt_0_143,.Wgt_0_144,.Wgt_0_145,.Wgt_0_146,.Wgt_0_147,.Wgt_0_148,.Wgt_0_149,.Wgt_0_150,.Wgt_0_151,.Wgt_0_152,.Wgt_0_153,.Wgt_0_154,.Wgt_0_155,.Wgt_0_156,.Wgt_0_157,.Wgt_0_158,.Wgt_0_159,.Wgt_0_160,.Wgt_0_161,.Wgt_0_162,.Wgt_0_163,.Wgt_0_164,.Wgt_0_165,.Wgt_0_166,.Wgt_0_167,.Wgt_0_168,.Wgt_0_169,.Wgt_0_170,.Wgt_0_171,.Wgt_0_172,.Wgt_0_173,.Wgt_0_174,.Wgt_0_175,.Wgt_0_176,.Wgt_0_177,.Wgt_0_178,.Wgt_0_179,.Wgt_0_180,.Wgt_0_181,.Wgt_0_182,.Wgt_0_183,.Wgt_0_184,.Wgt_0_185,.Wgt_0_186,.Wgt_0_187,.Wgt_0_188,.Wgt_0_189,.Wgt_0_190,.Wgt_0_191,.Wgt_0_192,.Wgt_0_193,.Wgt_0_194,.Wgt_0_195,.Wgt_0_196,.Wgt_0_197,.Wgt_0_198,.Wgt_0_199,.Wgt_0_200,.Wgt_0_201,.Wgt_0_202,.Wgt_0_203,.Wgt_0_204,.Wgt_0_205,.Wgt_0_206,.Wgt_0_207,.Wgt_0_208,.Wgt_0_209,.Wgt_0_210,.Wgt_0_211,.Wgt_0_212,.Wgt_0_213,.Wgt_0_214,.Wgt_0_215,.Wgt_0_216,.Wgt_0_217,.Wgt_0_218,.Wgt_0_219,.Wgt_0_220,.Wgt_0_221,.Wgt_0_222,.Wgt_0_223,.Wgt_0_224,.Wgt_0_225,.Wgt_0_226,.Wgt_0_227,.Wgt_0_228,.Wgt_0_229,.Wgt_0_230,.Wgt_0_231,.Wgt_0_232,.Wgt_0_233,.Wgt_0_234,.Wgt_0_235,.Wgt_0_236,.Wgt_0_237,.Wgt_0_238,.Wgt_0_239,.Wgt_0_240,.Wgt_0_241,.Wgt_0_242,.Wgt_0_243,.Wgt_0_244,.Wgt_0_245,.Wgt_0_246,.Wgt_0_247,.Wgt_0_248,.Wgt_0_249,.Wgt_0_250,.Wgt_0_251,.Wgt_0_252,.Wgt_0_253,.Wgt_0_254,.Wgt_0_255,.Wgt_0_256,.Wgt_0_257,.Wgt_0_258,.Wgt_0_259,.Wgt_0_260,.Wgt_0_261,.Wgt_0_262,.Wgt_0_263,.Wgt_0_264,.Wgt_0_265,.Wgt_0_266,.Wgt_0_267,.Wgt_0_268,.Wgt_0_269,.Wgt_0_270,.Wgt_0_271,.Wgt_0_272,.Wgt_0_273,.Wgt_0_274,.Wgt_0_275,.Wgt_0_276,.Wgt_0_277,.Wgt_0_278,.Wgt_0_279,.Wgt_0_280,.Wgt_0_281,.Wgt_0_282,.Wgt_0_283,.Wgt_0_284,.Wgt_0_285,.Wgt_0_286,.Wgt_0_287,.Wgt_0_288,.Wgt_0_289,.Wgt_0_290,.Wgt_0_291,.Wgt_0_292,.Wgt_0_293,.Wgt_0_294,.Wgt_0_295,.Wgt_0_296,.Wgt_0_297,.Wgt_0_298,.Wgt_0_299,.Wgt_0_300,.Wgt_0_301,.Wgt_0_302,.Wgt_0_303,.Wgt_0_304,.Wgt_0_305,.Wgt_0_306,.Wgt_0_307,.Wgt_0_308,.Wgt_0_309,.Wgt_0_310,.Wgt_0_311,.Wgt_0_312,.Wgt_0_313,.Wgt_0_314,.Wgt_0_315,.Wgt_0_316,.Wgt_0_317,.Wgt_0_318,.Wgt_0_319,.Wgt_0_320,.Wgt_0_321,.Wgt_0_322,.Wgt_0_323,.Wgt_0_324,.Wgt_0_325,.Wgt_0_326,.Wgt_0_327,.Wgt_0_328,.Wgt_0_329,.Wgt_0_330,.Wgt_0_331,.Wgt_0_332,.Wgt_0_333,.Wgt_0_334,.Wgt_0_335,.Wgt_0_336,.Wgt_0_337,.Wgt_0_338,.Wgt_0_339,.Wgt_0_340,.Wgt_0_341,.Wgt_0_342,.Wgt_0_343,.Wgt_0_344,.Wgt_0_345,.Wgt_0_346,.Wgt_0_347,.Wgt_0_348,.Wgt_0_349,.Wgt_0_350,.Wgt_0_351,.Wgt_0_352,.Wgt_0_353,.Wgt_0_354,.Wgt_0_355,.Wgt_0_356,.Wgt_0_357,.Wgt_0_358,.Wgt_0_359,.Wgt_0_360,.Wgt_0_361,.Wgt_0_362,.Wgt_0_363,.Wgt_0_364,.Wgt_0_365,.Wgt_0_366,.Wgt_0_367,.Wgt_0_368,.Wgt_0_369,.Wgt_0_370,.Wgt_0_371,.Wgt_0_372,.Wgt_0_373,.Wgt_0_374,.Wgt_0_375,.Wgt_0_376,.Wgt_0_377,.Wgt_0_378,.Wgt_0_379,.Wgt_0_380,.Wgt_0_381,.Wgt_0_382,.Wgt_0_383,.Wgt_0_384,.Wgt_0_385,.Wgt_0_386,.Wgt_0_387,.Wgt_0_388,.Wgt_0_389,.Wgt_0_390,.Wgt_0_391,.Wgt_0_392,.Wgt_0_393,.Wgt_0_394,.Wgt_0_395,.Wgt_0_396,.Wgt_0_397,.Wgt_0_398,.Wgt_0_399,.Wgt_0_400,.Wgt_0_401,.Wgt_0_402,.Wgt_0_403,.Wgt_0_404,.Wgt_0_405,.Wgt_0_406,.Wgt_0_407,.Wgt_0_408,.Wgt_0_409,.Wgt_0_410,.Wgt_0_411,.Wgt_0_412,.Wgt_0_413,.Wgt_0_414,.Wgt_0_415,.Wgt_0_416,.Wgt_0_417,.Wgt_0_418,.Wgt_0_419,.Wgt_0_420,.Wgt_0_421,.Wgt_0_422,.Wgt_0_423,.Wgt_0_424,.Wgt_0_425,.Wgt_0_426,.Wgt_0_427,.Wgt_0_428,.Wgt_0_429,.Wgt_0_430,.Wgt_0_431,.Wgt_0_432,.Wgt_0_433,.Wgt_0_434,.Wgt_0_435,.Wgt_0_436,.Wgt_0_437,.Wgt_0_438,.Wgt_0_439,.Wgt_0_440,.Wgt_0_441,.Wgt_0_442,.Wgt_0_443,.Wgt_0_444,.Wgt_0_445,.Wgt_0_446,.Wgt_0_447,.Wgt_0_448,.Wgt_0_449,.Wgt_0_450,.Wgt_0_451,.Wgt_0_452,.Wgt_0_453,.Wgt_0_454,.Wgt_0_455,.Wgt_0_456,.Wgt_0_457,.Wgt_0_458,.Wgt_0_459,.Wgt_0_460,.Wgt_0_461,.Wgt_0_462,.Wgt_0_463,.Wgt_0_464,.Wgt_0_465,.Wgt_0_466,.Wgt_0_467,.Wgt_0_468,.Wgt_0_469,.Wgt_0_470,.Wgt_0_471,.Wgt_0_472,.Wgt_0_473,.Wgt_0_474,.Wgt_0_475,.Wgt_0_476,.Wgt_0_477,.Wgt_0_478,.Wgt_0_479,.Wgt_0_480,.Wgt_0_481,.Wgt_0_482,.Wgt_0_483,.Wgt_0_484,.Wgt_0_485,.Wgt_0_486,.Wgt_0_487,.Wgt_0_488,.Wgt_0_489,.Wgt_0_490,.Wgt_0_491,.Wgt_0_492,.Wgt_0_493,.Wgt_0_494,.Wgt_0_495,.Wgt_0_496,.Wgt_0_497,.Wgt_0_498,.Wgt_0_499,.Wgt_0_500,.Wgt_0_501,.Wgt_0_502,.Wgt_0_503,.Wgt_0_504,.Wgt_0_505,.Wgt_0_506,.Wgt_0_507,.Wgt_0_508,.Wgt_0_509,.Wgt_0_510,.Wgt_0_511,.Wgt_0_512,.Wgt_0_513,.Wgt_0_514,.Wgt_0_515,.Wgt_0_516,.Wgt_0_517,.Wgt_0_518,.Wgt_0_519,.Wgt_0_520,.Wgt_0_521,.Wgt_0_522,.Wgt_0_523,.Wgt_0_524,.Wgt_0_525,.Wgt_0_526,.Wgt_0_527,.Wgt_0_528,.Wgt_0_529,.Wgt_0_530,.Wgt_0_531,.Wgt_0_532,.Wgt_0_533,.Wgt_0_534,.Wgt_0_535,.Wgt_0_536,.Wgt_0_537,.Wgt_0_538,.Wgt_0_539,.Wgt_0_540,.Wgt_0_541,.Wgt_0_542,.Wgt_0_543,.Wgt_0_544,.Wgt_0_545,.Wgt_0_546,.Wgt_0_547,.Wgt_0_548,.Wgt_0_549,.Wgt_0_550,.Wgt_0_551,.Wgt_0_552,.Wgt_0_553,.Wgt_0_554,.Wgt_0_555,.Wgt_0_556,.Wgt_0_557,.Wgt_0_558,.Wgt_0_559,.Wgt_0_560,.Wgt_0_561,.Wgt_0_562,.Wgt_0_563,.Wgt_0_564,.Wgt_0_565,.Wgt_0_566,.Wgt_0_567,.Wgt_0_568,.Wgt_0_569,.Wgt_0_570,.Wgt_0_571,.Wgt_0_572,.Wgt_0_573,.Wgt_0_574,.Wgt_0_575,.Wgt_0_576,.Wgt_0_577,.Wgt_0_578,.Wgt_0_579,.Wgt_0_580,.Wgt_0_581,.Wgt_0_582,.Wgt_0_583,.Wgt_0_584,.Wgt_0_585,.Wgt_0_586,.Wgt_0_587,.Wgt_0_588,.Wgt_0_589,.Wgt_0_590,.Wgt_0_591,.Wgt_0_592,.Wgt_0_593,.Wgt_0_594,.Wgt_0_595,.Wgt_0_596,.Wgt_0_597,.Wgt_0_598,.Wgt_0_599,.Wgt_0_600,.Wgt_0_601,.Wgt_0_602,.Wgt_0_603,.Wgt_0_604,.Wgt_0_605,.Wgt_0_606,.Wgt_0_607,.Wgt_0_608,.Wgt_0_609,.Wgt_0_610,.Wgt_0_611,.Wgt_0_612,.Wgt_0_613,.Wgt_0_614,.Wgt_0_615,.Wgt_0_616,.Wgt_0_617,.Wgt_0_618,.Wgt_0_619,.Wgt_0_620,.Wgt_0_621,.Wgt_0_622,.Wgt_0_623,.Wgt_0_624,.Wgt_0_625,.Wgt_0_626,.Wgt_0_627,.Wgt_0_628,.Wgt_0_629,.Wgt_0_630,.Wgt_0_631,.Wgt_0_632,.Wgt_0_633,.Wgt_0_634,.Wgt_0_635,.Wgt_0_636,.Wgt_0_637,.Wgt_0_638,.Wgt_0_639,.Wgt_0_640,.Wgt_0_641,.Wgt_0_642,.Wgt_0_643,.Wgt_0_644,.Wgt_0_645,.Wgt_0_646,.Wgt_0_647,.Wgt_0_648,.Wgt_0_649,.Wgt_0_650,.Wgt_0_651,.Wgt_0_652,.Wgt_0_653,.Wgt_0_654,.Wgt_0_655,.Wgt_0_656,.Wgt_0_657,.Wgt_0_658,.Wgt_0_659,.Wgt_0_660,.Wgt_0_661,.Wgt_0_662,.Wgt_0_663,.Wgt_0_664,.Wgt_0_665,.Wgt_0_666,.Wgt_0_667,.Wgt_0_668,.Wgt_0_669,.Wgt_0_670,.Wgt_0_671,.Wgt_0_672,.Wgt_0_673,.Wgt_0_674,.Wgt_0_675,.Wgt_0_676,.Wgt_0_677,.Wgt_0_678,.Wgt_0_679,.Wgt_0_680,.Wgt_0_681,.Wgt_0_682,.Wgt_0_683,.Wgt_0_684,.Wgt_0_685,.Wgt_0_686,.Wgt_0_687,.Wgt_0_688,.Wgt_0_689,.Wgt_0_690,.Wgt_0_691,.Wgt_0_692,.Wgt_0_693,.Wgt_0_694,.Wgt_0_695,.Wgt_0_696,.Wgt_0_697,.Wgt_0_698,.Wgt_0_699,.Wgt_0_700,.Wgt_0_701,.Wgt_0_702,.Wgt_0_703,.Wgt_0_704,.Wgt_0_705,.Wgt_0_706,.Wgt_0_707,.Wgt_0_708,.Wgt_0_709,.Wgt_0_710,.Wgt_0_711,.Wgt_0_712,.Wgt_0_713,.Wgt_0_714,.Wgt_0_715,.Wgt_0_716,.Wgt_0_717,.Wgt_0_718,.Wgt_0_719,.Wgt_0_720,.Wgt_0_721,.Wgt_0_722,.Wgt_0_723,.Wgt_0_724,.Wgt_0_725,.Wgt_0_726,.Wgt_0_727,.Wgt_0_728,.Wgt_0_729,.Wgt_0_730,.Wgt_0_731,.Wgt_0_732,.Wgt_0_733,.Wgt_0_734,.Wgt_0_735,.Wgt_0_736,.Wgt_0_737,.Wgt_0_738,.Wgt_0_739,.Wgt_0_740,.Wgt_0_741,.Wgt_0_742,.Wgt_0_743,.Wgt_0_744,.Wgt_0_745,.Wgt_0_746,.Wgt_0_747,.Wgt_0_748,.Wgt_0_749,.Wgt_0_750,.Wgt_0_751,.Wgt_0_752,.Wgt_0_753,.Wgt_0_754,.Wgt_0_755,.Wgt_0_756,.Wgt_0_757,.Wgt_0_758,.Wgt_0_759,.Wgt_0_760,.Wgt_0_761,.Wgt_0_762,.Wgt_0_763,.Wgt_0_764,.Wgt_0_765,.Wgt_0_766,.Wgt_0_767,.Wgt_0_768,.Wgt_0_769,.Wgt_0_770,.Wgt_0_771,.Wgt_0_772,.Wgt_0_773,.Wgt_0_774,.Wgt_0_775,.Wgt_0_776,.Wgt_0_777,.Wgt_0_778,.Wgt_0_779,.Wgt_0_780,.Wgt_0_781,.Wgt_0_782,.Wgt_0_783,.Wgt_0_784,
.Wgt_1_0,.Wgt_1_1,.Wgt_1_2,.Wgt_1_3,.Wgt_1_4,.Wgt_1_5,.Wgt_1_6,.Wgt_1_7,.Wgt_1_8,.Wgt_1_9,.Wgt_1_10,.Wgt_1_11,.Wgt_1_12,.Wgt_1_13,.Wgt_1_14,.Wgt_1_15,.Wgt_1_16,.Wgt_1_17,.Wgt_1_18,.Wgt_1_19,.Wgt_1_20,.Wgt_1_21,.Wgt_1_22,.Wgt_1_23,.Wgt_1_24,.Wgt_1_25,.Wgt_1_26,.Wgt_1_27,.Wgt_1_28,.Wgt_1_29,.Wgt_1_30,.Wgt_1_31,.Wgt_1_32,.Wgt_1_33,.Wgt_1_34,.Wgt_1_35,.Wgt_1_36,.Wgt_1_37,.Wgt_1_38,.Wgt_1_39,.Wgt_1_40,.Wgt_1_41,.Wgt_1_42,.Wgt_1_43,.Wgt_1_44,.Wgt_1_45,.Wgt_1_46,.Wgt_1_47,.Wgt_1_48,.Wgt_1_49,.Wgt_1_50,.Wgt_1_51,.Wgt_1_52,.Wgt_1_53,.Wgt_1_54,.Wgt_1_55,.Wgt_1_56,.Wgt_1_57,.Wgt_1_58,.Wgt_1_59,.Wgt_1_60,.Wgt_1_61,.Wgt_1_62,.Wgt_1_63,.Wgt_1_64,.Wgt_1_65,.Wgt_1_66,.Wgt_1_67,.Wgt_1_68,.Wgt_1_69,.Wgt_1_70,.Wgt_1_71,.Wgt_1_72,.Wgt_1_73,.Wgt_1_74,.Wgt_1_75,.Wgt_1_76,.Wgt_1_77,.Wgt_1_78,.Wgt_1_79,.Wgt_1_80,.Wgt_1_81,.Wgt_1_82,.Wgt_1_83,.Wgt_1_84,.Wgt_1_85,.Wgt_1_86,.Wgt_1_87,.Wgt_1_88,.Wgt_1_89,.Wgt_1_90,.Wgt_1_91,.Wgt_1_92,.Wgt_1_93,.Wgt_1_94,.Wgt_1_95,.Wgt_1_96,.Wgt_1_97,.Wgt_1_98,.Wgt_1_99,.Wgt_1_100,.Wgt_1_101,.Wgt_1_102,.Wgt_1_103,.Wgt_1_104,.Wgt_1_105,.Wgt_1_106,.Wgt_1_107,.Wgt_1_108,.Wgt_1_109,.Wgt_1_110,.Wgt_1_111,.Wgt_1_112,.Wgt_1_113,.Wgt_1_114,.Wgt_1_115,.Wgt_1_116,.Wgt_1_117,.Wgt_1_118,.Wgt_1_119,.Wgt_1_120,.Wgt_1_121,.Wgt_1_122,.Wgt_1_123,.Wgt_1_124,.Wgt_1_125,.Wgt_1_126,.Wgt_1_127,.Wgt_1_128,.Wgt_1_129,.Wgt_1_130,.Wgt_1_131,.Wgt_1_132,.Wgt_1_133,.Wgt_1_134,.Wgt_1_135,.Wgt_1_136,.Wgt_1_137,.Wgt_1_138,.Wgt_1_139,.Wgt_1_140,.Wgt_1_141,.Wgt_1_142,.Wgt_1_143,.Wgt_1_144,.Wgt_1_145,.Wgt_1_146,.Wgt_1_147,.Wgt_1_148,.Wgt_1_149,.Wgt_1_150,.Wgt_1_151,.Wgt_1_152,.Wgt_1_153,.Wgt_1_154,.Wgt_1_155,.Wgt_1_156,.Wgt_1_157,.Wgt_1_158,.Wgt_1_159,.Wgt_1_160,.Wgt_1_161,.Wgt_1_162,.Wgt_1_163,.Wgt_1_164,.Wgt_1_165,.Wgt_1_166,.Wgt_1_167,.Wgt_1_168,.Wgt_1_169,.Wgt_1_170,.Wgt_1_171,.Wgt_1_172,.Wgt_1_173,.Wgt_1_174,.Wgt_1_175,.Wgt_1_176,.Wgt_1_177,.Wgt_1_178,.Wgt_1_179,.Wgt_1_180,.Wgt_1_181,.Wgt_1_182,.Wgt_1_183,.Wgt_1_184,.Wgt_1_185,.Wgt_1_186,.Wgt_1_187,.Wgt_1_188,.Wgt_1_189,.Wgt_1_190,.Wgt_1_191,.Wgt_1_192,.Wgt_1_193,.Wgt_1_194,.Wgt_1_195,.Wgt_1_196,.Wgt_1_197,.Wgt_1_198,.Wgt_1_199,.Wgt_1_200,.Wgt_1_201,.Wgt_1_202,.Wgt_1_203,.Wgt_1_204,.Wgt_1_205,.Wgt_1_206,.Wgt_1_207,.Wgt_1_208,.Wgt_1_209,.Wgt_1_210,.Wgt_1_211,.Wgt_1_212,.Wgt_1_213,.Wgt_1_214,.Wgt_1_215,.Wgt_1_216,.Wgt_1_217,.Wgt_1_218,.Wgt_1_219,.Wgt_1_220,.Wgt_1_221,.Wgt_1_222,.Wgt_1_223,.Wgt_1_224,.Wgt_1_225,.Wgt_1_226,.Wgt_1_227,.Wgt_1_228,.Wgt_1_229,.Wgt_1_230,.Wgt_1_231,.Wgt_1_232,.Wgt_1_233,.Wgt_1_234,.Wgt_1_235,.Wgt_1_236,.Wgt_1_237,.Wgt_1_238,.Wgt_1_239,.Wgt_1_240,.Wgt_1_241,.Wgt_1_242,.Wgt_1_243,.Wgt_1_244,.Wgt_1_245,.Wgt_1_246,.Wgt_1_247,.Wgt_1_248,.Wgt_1_249,.Wgt_1_250,.Wgt_1_251,.Wgt_1_252,.Wgt_1_253,.Wgt_1_254,.Wgt_1_255,.Wgt_1_256,.Wgt_1_257,.Wgt_1_258,.Wgt_1_259,.Wgt_1_260,.Wgt_1_261,.Wgt_1_262,.Wgt_1_263,.Wgt_1_264,.Wgt_1_265,.Wgt_1_266,.Wgt_1_267,.Wgt_1_268,.Wgt_1_269,.Wgt_1_270,.Wgt_1_271,.Wgt_1_272,.Wgt_1_273,.Wgt_1_274,.Wgt_1_275,.Wgt_1_276,.Wgt_1_277,.Wgt_1_278,.Wgt_1_279,.Wgt_1_280,.Wgt_1_281,.Wgt_1_282,.Wgt_1_283,.Wgt_1_284,.Wgt_1_285,.Wgt_1_286,.Wgt_1_287,.Wgt_1_288,.Wgt_1_289,.Wgt_1_290,.Wgt_1_291,.Wgt_1_292,.Wgt_1_293,.Wgt_1_294,.Wgt_1_295,.Wgt_1_296,.Wgt_1_297,.Wgt_1_298,.Wgt_1_299,.Wgt_1_300,.Wgt_1_301,.Wgt_1_302,.Wgt_1_303,.Wgt_1_304,.Wgt_1_305,.Wgt_1_306,.Wgt_1_307,.Wgt_1_308,.Wgt_1_309,.Wgt_1_310,.Wgt_1_311,.Wgt_1_312,.Wgt_1_313,.Wgt_1_314,.Wgt_1_315,.Wgt_1_316,.Wgt_1_317,.Wgt_1_318,.Wgt_1_319,.Wgt_1_320,.Wgt_1_321,.Wgt_1_322,.Wgt_1_323,.Wgt_1_324,.Wgt_1_325,.Wgt_1_326,.Wgt_1_327,.Wgt_1_328,.Wgt_1_329,.Wgt_1_330,.Wgt_1_331,.Wgt_1_332,.Wgt_1_333,.Wgt_1_334,.Wgt_1_335,.Wgt_1_336,.Wgt_1_337,.Wgt_1_338,.Wgt_1_339,.Wgt_1_340,.Wgt_1_341,.Wgt_1_342,.Wgt_1_343,.Wgt_1_344,.Wgt_1_345,.Wgt_1_346,.Wgt_1_347,.Wgt_1_348,.Wgt_1_349,.Wgt_1_350,.Wgt_1_351,.Wgt_1_352,.Wgt_1_353,.Wgt_1_354,.Wgt_1_355,.Wgt_1_356,.Wgt_1_357,.Wgt_1_358,.Wgt_1_359,.Wgt_1_360,.Wgt_1_361,.Wgt_1_362,.Wgt_1_363,.Wgt_1_364,.Wgt_1_365,.Wgt_1_366,.Wgt_1_367,.Wgt_1_368,.Wgt_1_369,.Wgt_1_370,.Wgt_1_371,.Wgt_1_372,.Wgt_1_373,.Wgt_1_374,.Wgt_1_375,.Wgt_1_376,.Wgt_1_377,.Wgt_1_378,.Wgt_1_379,.Wgt_1_380,.Wgt_1_381,.Wgt_1_382,.Wgt_1_383,.Wgt_1_384,.Wgt_1_385,.Wgt_1_386,.Wgt_1_387,.Wgt_1_388,.Wgt_1_389,.Wgt_1_390,.Wgt_1_391,.Wgt_1_392,.Wgt_1_393,.Wgt_1_394,.Wgt_1_395,.Wgt_1_396,.Wgt_1_397,.Wgt_1_398,.Wgt_1_399,.Wgt_1_400,.Wgt_1_401,.Wgt_1_402,.Wgt_1_403,.Wgt_1_404,.Wgt_1_405,.Wgt_1_406,.Wgt_1_407,.Wgt_1_408,.Wgt_1_409,.Wgt_1_410,.Wgt_1_411,.Wgt_1_412,.Wgt_1_413,.Wgt_1_414,.Wgt_1_415,.Wgt_1_416,.Wgt_1_417,.Wgt_1_418,.Wgt_1_419,.Wgt_1_420,.Wgt_1_421,.Wgt_1_422,.Wgt_1_423,.Wgt_1_424,.Wgt_1_425,.Wgt_1_426,.Wgt_1_427,.Wgt_1_428,.Wgt_1_429,.Wgt_1_430,.Wgt_1_431,.Wgt_1_432,.Wgt_1_433,.Wgt_1_434,.Wgt_1_435,.Wgt_1_436,.Wgt_1_437,.Wgt_1_438,.Wgt_1_439,.Wgt_1_440,.Wgt_1_441,.Wgt_1_442,.Wgt_1_443,.Wgt_1_444,.Wgt_1_445,.Wgt_1_446,.Wgt_1_447,.Wgt_1_448,.Wgt_1_449,.Wgt_1_450,.Wgt_1_451,.Wgt_1_452,.Wgt_1_453,.Wgt_1_454,.Wgt_1_455,.Wgt_1_456,.Wgt_1_457,.Wgt_1_458,.Wgt_1_459,.Wgt_1_460,.Wgt_1_461,.Wgt_1_462,.Wgt_1_463,.Wgt_1_464,.Wgt_1_465,.Wgt_1_466,.Wgt_1_467,.Wgt_1_468,.Wgt_1_469,.Wgt_1_470,.Wgt_1_471,.Wgt_1_472,.Wgt_1_473,.Wgt_1_474,.Wgt_1_475,.Wgt_1_476,.Wgt_1_477,.Wgt_1_478,.Wgt_1_479,.Wgt_1_480,.Wgt_1_481,.Wgt_1_482,.Wgt_1_483,.Wgt_1_484,.Wgt_1_485,.Wgt_1_486,.Wgt_1_487,.Wgt_1_488,.Wgt_1_489,.Wgt_1_490,.Wgt_1_491,.Wgt_1_492,.Wgt_1_493,.Wgt_1_494,.Wgt_1_495,.Wgt_1_496,.Wgt_1_497,.Wgt_1_498,.Wgt_1_499,.Wgt_1_500,.Wgt_1_501,.Wgt_1_502,.Wgt_1_503,.Wgt_1_504,.Wgt_1_505,.Wgt_1_506,.Wgt_1_507,.Wgt_1_508,.Wgt_1_509,.Wgt_1_510,.Wgt_1_511,.Wgt_1_512,.Wgt_1_513,.Wgt_1_514,.Wgt_1_515,.Wgt_1_516,.Wgt_1_517,.Wgt_1_518,.Wgt_1_519,.Wgt_1_520,.Wgt_1_521,.Wgt_1_522,.Wgt_1_523,.Wgt_1_524,.Wgt_1_525,.Wgt_1_526,.Wgt_1_527,.Wgt_1_528,.Wgt_1_529,.Wgt_1_530,.Wgt_1_531,.Wgt_1_532,.Wgt_1_533,.Wgt_1_534,.Wgt_1_535,.Wgt_1_536,.Wgt_1_537,.Wgt_1_538,.Wgt_1_539,.Wgt_1_540,.Wgt_1_541,.Wgt_1_542,.Wgt_1_543,.Wgt_1_544,.Wgt_1_545,.Wgt_1_546,.Wgt_1_547,.Wgt_1_548,.Wgt_1_549,.Wgt_1_550,.Wgt_1_551,.Wgt_1_552,.Wgt_1_553,.Wgt_1_554,.Wgt_1_555,.Wgt_1_556,.Wgt_1_557,.Wgt_1_558,.Wgt_1_559,.Wgt_1_560,.Wgt_1_561,.Wgt_1_562,.Wgt_1_563,.Wgt_1_564,.Wgt_1_565,.Wgt_1_566,.Wgt_1_567,.Wgt_1_568,.Wgt_1_569,.Wgt_1_570,.Wgt_1_571,.Wgt_1_572,.Wgt_1_573,.Wgt_1_574,.Wgt_1_575,.Wgt_1_576,.Wgt_1_577,.Wgt_1_578,.Wgt_1_579,.Wgt_1_580,.Wgt_1_581,.Wgt_1_582,.Wgt_1_583,.Wgt_1_584,.Wgt_1_585,.Wgt_1_586,.Wgt_1_587,.Wgt_1_588,.Wgt_1_589,.Wgt_1_590,.Wgt_1_591,.Wgt_1_592,.Wgt_1_593,.Wgt_1_594,.Wgt_1_595,.Wgt_1_596,.Wgt_1_597,.Wgt_1_598,.Wgt_1_599,.Wgt_1_600,.Wgt_1_601,.Wgt_1_602,.Wgt_1_603,.Wgt_1_604,.Wgt_1_605,.Wgt_1_606,.Wgt_1_607,.Wgt_1_608,.Wgt_1_609,.Wgt_1_610,.Wgt_1_611,.Wgt_1_612,.Wgt_1_613,.Wgt_1_614,.Wgt_1_615,.Wgt_1_616,.Wgt_1_617,.Wgt_1_618,.Wgt_1_619,.Wgt_1_620,.Wgt_1_621,.Wgt_1_622,.Wgt_1_623,.Wgt_1_624,.Wgt_1_625,.Wgt_1_626,.Wgt_1_627,.Wgt_1_628,.Wgt_1_629,.Wgt_1_630,.Wgt_1_631,.Wgt_1_632,.Wgt_1_633,.Wgt_1_634,.Wgt_1_635,.Wgt_1_636,.Wgt_1_637,.Wgt_1_638,.Wgt_1_639,.Wgt_1_640,.Wgt_1_641,.Wgt_1_642,.Wgt_1_643,.Wgt_1_644,.Wgt_1_645,.Wgt_1_646,.Wgt_1_647,.Wgt_1_648,.Wgt_1_649,.Wgt_1_650,.Wgt_1_651,.Wgt_1_652,.Wgt_1_653,.Wgt_1_654,.Wgt_1_655,.Wgt_1_656,.Wgt_1_657,.Wgt_1_658,.Wgt_1_659,.Wgt_1_660,.Wgt_1_661,.Wgt_1_662,.Wgt_1_663,.Wgt_1_664,.Wgt_1_665,.Wgt_1_666,.Wgt_1_667,.Wgt_1_668,.Wgt_1_669,.Wgt_1_670,.Wgt_1_671,.Wgt_1_672,.Wgt_1_673,.Wgt_1_674,.Wgt_1_675,.Wgt_1_676,.Wgt_1_677,.Wgt_1_678,.Wgt_1_679,.Wgt_1_680,.Wgt_1_681,.Wgt_1_682,.Wgt_1_683,.Wgt_1_684,.Wgt_1_685,.Wgt_1_686,.Wgt_1_687,.Wgt_1_688,.Wgt_1_689,.Wgt_1_690,.Wgt_1_691,.Wgt_1_692,.Wgt_1_693,.Wgt_1_694,.Wgt_1_695,.Wgt_1_696,.Wgt_1_697,.Wgt_1_698,.Wgt_1_699,.Wgt_1_700,.Wgt_1_701,.Wgt_1_702,.Wgt_1_703,.Wgt_1_704,.Wgt_1_705,.Wgt_1_706,.Wgt_1_707,.Wgt_1_708,.Wgt_1_709,.Wgt_1_710,.Wgt_1_711,.Wgt_1_712,.Wgt_1_713,.Wgt_1_714,.Wgt_1_715,.Wgt_1_716,.Wgt_1_717,.Wgt_1_718,.Wgt_1_719,.Wgt_1_720,.Wgt_1_721,.Wgt_1_722,.Wgt_1_723,.Wgt_1_724,.Wgt_1_725,.Wgt_1_726,.Wgt_1_727,.Wgt_1_728,.Wgt_1_729,.Wgt_1_730,.Wgt_1_731,.Wgt_1_732,.Wgt_1_733,.Wgt_1_734,.Wgt_1_735,.Wgt_1_736,.Wgt_1_737,.Wgt_1_738,.Wgt_1_739,.Wgt_1_740,.Wgt_1_741,.Wgt_1_742,.Wgt_1_743,.Wgt_1_744,.Wgt_1_745,.Wgt_1_746,.Wgt_1_747,.Wgt_1_748,.Wgt_1_749,.Wgt_1_750,.Wgt_1_751,.Wgt_1_752,.Wgt_1_753,.Wgt_1_754,.Wgt_1_755,.Wgt_1_756,.Wgt_1_757,.Wgt_1_758,.Wgt_1_759,.Wgt_1_760,.Wgt_1_761,.Wgt_1_762,.Wgt_1_763,.Wgt_1_764,.Wgt_1_765,.Wgt_1_766,.Wgt_1_767,.Wgt_1_768,.Wgt_1_769,.Wgt_1_770,.Wgt_1_771,.Wgt_1_772,.Wgt_1_773,.Wgt_1_774,.Wgt_1_775,.Wgt_1_776,.Wgt_1_777,.Wgt_1_778,.Wgt_1_779,.Wgt_1_780,.Wgt_1_781,.Wgt_1_782,.Wgt_1_783,.Wgt_1_784,
.Wgt_2_0,.Wgt_2_1,.Wgt_2_2,.Wgt_2_3,.Wgt_2_4,.Wgt_2_5,.Wgt_2_6,.Wgt_2_7,.Wgt_2_8,.Wgt_2_9,.Wgt_2_10,.Wgt_2_11,.Wgt_2_12,.Wgt_2_13,.Wgt_2_14,.Wgt_2_15,.Wgt_2_16,.Wgt_2_17,.Wgt_2_18,.Wgt_2_19,.Wgt_2_20,.Wgt_2_21,.Wgt_2_22,.Wgt_2_23,.Wgt_2_24,.Wgt_2_25,.Wgt_2_26,.Wgt_2_27,.Wgt_2_28,.Wgt_2_29,.Wgt_2_30,.Wgt_2_31,.Wgt_2_32,.Wgt_2_33,.Wgt_2_34,.Wgt_2_35,.Wgt_2_36,.Wgt_2_37,.Wgt_2_38,.Wgt_2_39,.Wgt_2_40,.Wgt_2_41,.Wgt_2_42,.Wgt_2_43,.Wgt_2_44,.Wgt_2_45,.Wgt_2_46,.Wgt_2_47,.Wgt_2_48,.Wgt_2_49,.Wgt_2_50,.Wgt_2_51,.Wgt_2_52,.Wgt_2_53,.Wgt_2_54,.Wgt_2_55,.Wgt_2_56,.Wgt_2_57,.Wgt_2_58,.Wgt_2_59,.Wgt_2_60,.Wgt_2_61,.Wgt_2_62,.Wgt_2_63,.Wgt_2_64,.Wgt_2_65,.Wgt_2_66,.Wgt_2_67,.Wgt_2_68,.Wgt_2_69,.Wgt_2_70,.Wgt_2_71,.Wgt_2_72,.Wgt_2_73,.Wgt_2_74,.Wgt_2_75,.Wgt_2_76,.Wgt_2_77,.Wgt_2_78,.Wgt_2_79,.Wgt_2_80,.Wgt_2_81,.Wgt_2_82,.Wgt_2_83,.Wgt_2_84,.Wgt_2_85,.Wgt_2_86,.Wgt_2_87,.Wgt_2_88,.Wgt_2_89,.Wgt_2_90,.Wgt_2_91,.Wgt_2_92,.Wgt_2_93,.Wgt_2_94,.Wgt_2_95,.Wgt_2_96,.Wgt_2_97,.Wgt_2_98,.Wgt_2_99,.Wgt_2_100,.Wgt_2_101,.Wgt_2_102,.Wgt_2_103,.Wgt_2_104,.Wgt_2_105,.Wgt_2_106,.Wgt_2_107,.Wgt_2_108,.Wgt_2_109,.Wgt_2_110,.Wgt_2_111,.Wgt_2_112,.Wgt_2_113,.Wgt_2_114,.Wgt_2_115,.Wgt_2_116,.Wgt_2_117,.Wgt_2_118,.Wgt_2_119,.Wgt_2_120,.Wgt_2_121,.Wgt_2_122,.Wgt_2_123,.Wgt_2_124,.Wgt_2_125,.Wgt_2_126,.Wgt_2_127,.Wgt_2_128,.Wgt_2_129,.Wgt_2_130,.Wgt_2_131,.Wgt_2_132,.Wgt_2_133,.Wgt_2_134,.Wgt_2_135,.Wgt_2_136,.Wgt_2_137,.Wgt_2_138,.Wgt_2_139,.Wgt_2_140,.Wgt_2_141,.Wgt_2_142,.Wgt_2_143,.Wgt_2_144,.Wgt_2_145,.Wgt_2_146,.Wgt_2_147,.Wgt_2_148,.Wgt_2_149,.Wgt_2_150,.Wgt_2_151,.Wgt_2_152,.Wgt_2_153,.Wgt_2_154,.Wgt_2_155,.Wgt_2_156,.Wgt_2_157,.Wgt_2_158,.Wgt_2_159,.Wgt_2_160,.Wgt_2_161,.Wgt_2_162,.Wgt_2_163,.Wgt_2_164,.Wgt_2_165,.Wgt_2_166,.Wgt_2_167,.Wgt_2_168,.Wgt_2_169,.Wgt_2_170,.Wgt_2_171,.Wgt_2_172,.Wgt_2_173,.Wgt_2_174,.Wgt_2_175,.Wgt_2_176,.Wgt_2_177,.Wgt_2_178,.Wgt_2_179,.Wgt_2_180,.Wgt_2_181,.Wgt_2_182,.Wgt_2_183,.Wgt_2_184,.Wgt_2_185,.Wgt_2_186,.Wgt_2_187,.Wgt_2_188,.Wgt_2_189,.Wgt_2_190,.Wgt_2_191,.Wgt_2_192,.Wgt_2_193,.Wgt_2_194,.Wgt_2_195,.Wgt_2_196,.Wgt_2_197,.Wgt_2_198,.Wgt_2_199,.Wgt_2_200,.Wgt_2_201,.Wgt_2_202,.Wgt_2_203,.Wgt_2_204,.Wgt_2_205,.Wgt_2_206,.Wgt_2_207,.Wgt_2_208,.Wgt_2_209,.Wgt_2_210,.Wgt_2_211,.Wgt_2_212,.Wgt_2_213,.Wgt_2_214,.Wgt_2_215,.Wgt_2_216,.Wgt_2_217,.Wgt_2_218,.Wgt_2_219,.Wgt_2_220,.Wgt_2_221,.Wgt_2_222,.Wgt_2_223,.Wgt_2_224,.Wgt_2_225,.Wgt_2_226,.Wgt_2_227,.Wgt_2_228,.Wgt_2_229,.Wgt_2_230,.Wgt_2_231,.Wgt_2_232,.Wgt_2_233,.Wgt_2_234,.Wgt_2_235,.Wgt_2_236,.Wgt_2_237,.Wgt_2_238,.Wgt_2_239,.Wgt_2_240,.Wgt_2_241,.Wgt_2_242,.Wgt_2_243,.Wgt_2_244,.Wgt_2_245,.Wgt_2_246,.Wgt_2_247,.Wgt_2_248,.Wgt_2_249,.Wgt_2_250,.Wgt_2_251,.Wgt_2_252,.Wgt_2_253,.Wgt_2_254,.Wgt_2_255,.Wgt_2_256,.Wgt_2_257,.Wgt_2_258,.Wgt_2_259,.Wgt_2_260,.Wgt_2_261,.Wgt_2_262,.Wgt_2_263,.Wgt_2_264,.Wgt_2_265,.Wgt_2_266,.Wgt_2_267,.Wgt_2_268,.Wgt_2_269,.Wgt_2_270,.Wgt_2_271,.Wgt_2_272,.Wgt_2_273,.Wgt_2_274,.Wgt_2_275,.Wgt_2_276,.Wgt_2_277,.Wgt_2_278,.Wgt_2_279,.Wgt_2_280,.Wgt_2_281,.Wgt_2_282,.Wgt_2_283,.Wgt_2_284,.Wgt_2_285,.Wgt_2_286,.Wgt_2_287,.Wgt_2_288,.Wgt_2_289,.Wgt_2_290,.Wgt_2_291,.Wgt_2_292,.Wgt_2_293,.Wgt_2_294,.Wgt_2_295,.Wgt_2_296,.Wgt_2_297,.Wgt_2_298,.Wgt_2_299,.Wgt_2_300,.Wgt_2_301,.Wgt_2_302,.Wgt_2_303,.Wgt_2_304,.Wgt_2_305,.Wgt_2_306,.Wgt_2_307,.Wgt_2_308,.Wgt_2_309,.Wgt_2_310,.Wgt_2_311,.Wgt_2_312,.Wgt_2_313,.Wgt_2_314,.Wgt_2_315,.Wgt_2_316,.Wgt_2_317,.Wgt_2_318,.Wgt_2_319,.Wgt_2_320,.Wgt_2_321,.Wgt_2_322,.Wgt_2_323,.Wgt_2_324,.Wgt_2_325,.Wgt_2_326,.Wgt_2_327,.Wgt_2_328,.Wgt_2_329,.Wgt_2_330,.Wgt_2_331,.Wgt_2_332,.Wgt_2_333,.Wgt_2_334,.Wgt_2_335,.Wgt_2_336,.Wgt_2_337,.Wgt_2_338,.Wgt_2_339,.Wgt_2_340,.Wgt_2_341,.Wgt_2_342,.Wgt_2_343,.Wgt_2_344,.Wgt_2_345,.Wgt_2_346,.Wgt_2_347,.Wgt_2_348,.Wgt_2_349,.Wgt_2_350,.Wgt_2_351,.Wgt_2_352,.Wgt_2_353,.Wgt_2_354,.Wgt_2_355,.Wgt_2_356,.Wgt_2_357,.Wgt_2_358,.Wgt_2_359,.Wgt_2_360,.Wgt_2_361,.Wgt_2_362,.Wgt_2_363,.Wgt_2_364,.Wgt_2_365,.Wgt_2_366,.Wgt_2_367,.Wgt_2_368,.Wgt_2_369,.Wgt_2_370,.Wgt_2_371,.Wgt_2_372,.Wgt_2_373,.Wgt_2_374,.Wgt_2_375,.Wgt_2_376,.Wgt_2_377,.Wgt_2_378,.Wgt_2_379,.Wgt_2_380,.Wgt_2_381,.Wgt_2_382,.Wgt_2_383,.Wgt_2_384,.Wgt_2_385,.Wgt_2_386,.Wgt_2_387,.Wgt_2_388,.Wgt_2_389,.Wgt_2_390,.Wgt_2_391,.Wgt_2_392,.Wgt_2_393,.Wgt_2_394,.Wgt_2_395,.Wgt_2_396,.Wgt_2_397,.Wgt_2_398,.Wgt_2_399,.Wgt_2_400,.Wgt_2_401,.Wgt_2_402,.Wgt_2_403,.Wgt_2_404,.Wgt_2_405,.Wgt_2_406,.Wgt_2_407,.Wgt_2_408,.Wgt_2_409,.Wgt_2_410,.Wgt_2_411,.Wgt_2_412,.Wgt_2_413,.Wgt_2_414,.Wgt_2_415,.Wgt_2_416,.Wgt_2_417,.Wgt_2_418,.Wgt_2_419,.Wgt_2_420,.Wgt_2_421,.Wgt_2_422,.Wgt_2_423,.Wgt_2_424,.Wgt_2_425,.Wgt_2_426,.Wgt_2_427,.Wgt_2_428,.Wgt_2_429,.Wgt_2_430,.Wgt_2_431,.Wgt_2_432,.Wgt_2_433,.Wgt_2_434,.Wgt_2_435,.Wgt_2_436,.Wgt_2_437,.Wgt_2_438,.Wgt_2_439,.Wgt_2_440,.Wgt_2_441,.Wgt_2_442,.Wgt_2_443,.Wgt_2_444,.Wgt_2_445,.Wgt_2_446,.Wgt_2_447,.Wgt_2_448,.Wgt_2_449,.Wgt_2_450,.Wgt_2_451,.Wgt_2_452,.Wgt_2_453,.Wgt_2_454,.Wgt_2_455,.Wgt_2_456,.Wgt_2_457,.Wgt_2_458,.Wgt_2_459,.Wgt_2_460,.Wgt_2_461,.Wgt_2_462,.Wgt_2_463,.Wgt_2_464,.Wgt_2_465,.Wgt_2_466,.Wgt_2_467,.Wgt_2_468,.Wgt_2_469,.Wgt_2_470,.Wgt_2_471,.Wgt_2_472,.Wgt_2_473,.Wgt_2_474,.Wgt_2_475,.Wgt_2_476,.Wgt_2_477,.Wgt_2_478,.Wgt_2_479,.Wgt_2_480,.Wgt_2_481,.Wgt_2_482,.Wgt_2_483,.Wgt_2_484,.Wgt_2_485,.Wgt_2_486,.Wgt_2_487,.Wgt_2_488,.Wgt_2_489,.Wgt_2_490,.Wgt_2_491,.Wgt_2_492,.Wgt_2_493,.Wgt_2_494,.Wgt_2_495,.Wgt_2_496,.Wgt_2_497,.Wgt_2_498,.Wgt_2_499,.Wgt_2_500,.Wgt_2_501,.Wgt_2_502,.Wgt_2_503,.Wgt_2_504,.Wgt_2_505,.Wgt_2_506,.Wgt_2_507,.Wgt_2_508,.Wgt_2_509,.Wgt_2_510,.Wgt_2_511,.Wgt_2_512,.Wgt_2_513,.Wgt_2_514,.Wgt_2_515,.Wgt_2_516,.Wgt_2_517,.Wgt_2_518,.Wgt_2_519,.Wgt_2_520,.Wgt_2_521,.Wgt_2_522,.Wgt_2_523,.Wgt_2_524,.Wgt_2_525,.Wgt_2_526,.Wgt_2_527,.Wgt_2_528,.Wgt_2_529,.Wgt_2_530,.Wgt_2_531,.Wgt_2_532,.Wgt_2_533,.Wgt_2_534,.Wgt_2_535,.Wgt_2_536,.Wgt_2_537,.Wgt_2_538,.Wgt_2_539,.Wgt_2_540,.Wgt_2_541,.Wgt_2_542,.Wgt_2_543,.Wgt_2_544,.Wgt_2_545,.Wgt_2_546,.Wgt_2_547,.Wgt_2_548,.Wgt_2_549,.Wgt_2_550,.Wgt_2_551,.Wgt_2_552,.Wgt_2_553,.Wgt_2_554,.Wgt_2_555,.Wgt_2_556,.Wgt_2_557,.Wgt_2_558,.Wgt_2_559,.Wgt_2_560,.Wgt_2_561,.Wgt_2_562,.Wgt_2_563,.Wgt_2_564,.Wgt_2_565,.Wgt_2_566,.Wgt_2_567,.Wgt_2_568,.Wgt_2_569,.Wgt_2_570,.Wgt_2_571,.Wgt_2_572,.Wgt_2_573,.Wgt_2_574,.Wgt_2_575,.Wgt_2_576,.Wgt_2_577,.Wgt_2_578,.Wgt_2_579,.Wgt_2_580,.Wgt_2_581,.Wgt_2_582,.Wgt_2_583,.Wgt_2_584,.Wgt_2_585,.Wgt_2_586,.Wgt_2_587,.Wgt_2_588,.Wgt_2_589,.Wgt_2_590,.Wgt_2_591,.Wgt_2_592,.Wgt_2_593,.Wgt_2_594,.Wgt_2_595,.Wgt_2_596,.Wgt_2_597,.Wgt_2_598,.Wgt_2_599,.Wgt_2_600,.Wgt_2_601,.Wgt_2_602,.Wgt_2_603,.Wgt_2_604,.Wgt_2_605,.Wgt_2_606,.Wgt_2_607,.Wgt_2_608,.Wgt_2_609,.Wgt_2_610,.Wgt_2_611,.Wgt_2_612,.Wgt_2_613,.Wgt_2_614,.Wgt_2_615,.Wgt_2_616,.Wgt_2_617,.Wgt_2_618,.Wgt_2_619,.Wgt_2_620,.Wgt_2_621,.Wgt_2_622,.Wgt_2_623,.Wgt_2_624,.Wgt_2_625,.Wgt_2_626,.Wgt_2_627,.Wgt_2_628,.Wgt_2_629,.Wgt_2_630,.Wgt_2_631,.Wgt_2_632,.Wgt_2_633,.Wgt_2_634,.Wgt_2_635,.Wgt_2_636,.Wgt_2_637,.Wgt_2_638,.Wgt_2_639,.Wgt_2_640,.Wgt_2_641,.Wgt_2_642,.Wgt_2_643,.Wgt_2_644,.Wgt_2_645,.Wgt_2_646,.Wgt_2_647,.Wgt_2_648,.Wgt_2_649,.Wgt_2_650,.Wgt_2_651,.Wgt_2_652,.Wgt_2_653,.Wgt_2_654,.Wgt_2_655,.Wgt_2_656,.Wgt_2_657,.Wgt_2_658,.Wgt_2_659,.Wgt_2_660,.Wgt_2_661,.Wgt_2_662,.Wgt_2_663,.Wgt_2_664,.Wgt_2_665,.Wgt_2_666,.Wgt_2_667,.Wgt_2_668,.Wgt_2_669,.Wgt_2_670,.Wgt_2_671,.Wgt_2_672,.Wgt_2_673,.Wgt_2_674,.Wgt_2_675,.Wgt_2_676,.Wgt_2_677,.Wgt_2_678,.Wgt_2_679,.Wgt_2_680,.Wgt_2_681,.Wgt_2_682,.Wgt_2_683,.Wgt_2_684,.Wgt_2_685,.Wgt_2_686,.Wgt_2_687,.Wgt_2_688,.Wgt_2_689,.Wgt_2_690,.Wgt_2_691,.Wgt_2_692,.Wgt_2_693,.Wgt_2_694,.Wgt_2_695,.Wgt_2_696,.Wgt_2_697,.Wgt_2_698,.Wgt_2_699,.Wgt_2_700,.Wgt_2_701,.Wgt_2_702,.Wgt_2_703,.Wgt_2_704,.Wgt_2_705,.Wgt_2_706,.Wgt_2_707,.Wgt_2_708,.Wgt_2_709,.Wgt_2_710,.Wgt_2_711,.Wgt_2_712,.Wgt_2_713,.Wgt_2_714,.Wgt_2_715,.Wgt_2_716,.Wgt_2_717,.Wgt_2_718,.Wgt_2_719,.Wgt_2_720,.Wgt_2_721,.Wgt_2_722,.Wgt_2_723,.Wgt_2_724,.Wgt_2_725,.Wgt_2_726,.Wgt_2_727,.Wgt_2_728,.Wgt_2_729,.Wgt_2_730,.Wgt_2_731,.Wgt_2_732,.Wgt_2_733,.Wgt_2_734,.Wgt_2_735,.Wgt_2_736,.Wgt_2_737,.Wgt_2_738,.Wgt_2_739,.Wgt_2_740,.Wgt_2_741,.Wgt_2_742,.Wgt_2_743,.Wgt_2_744,.Wgt_2_745,.Wgt_2_746,.Wgt_2_747,.Wgt_2_748,.Wgt_2_749,.Wgt_2_750,.Wgt_2_751,.Wgt_2_752,.Wgt_2_753,.Wgt_2_754,.Wgt_2_755,.Wgt_2_756,.Wgt_2_757,.Wgt_2_758,.Wgt_2_759,.Wgt_2_760,.Wgt_2_761,.Wgt_2_762,.Wgt_2_763,.Wgt_2_764,.Wgt_2_765,.Wgt_2_766,.Wgt_2_767,.Wgt_2_768,.Wgt_2_769,.Wgt_2_770,.Wgt_2_771,.Wgt_2_772,.Wgt_2_773,.Wgt_2_774,.Wgt_2_775,.Wgt_2_776,.Wgt_2_777,.Wgt_2_778,.Wgt_2_779,.Wgt_2_780,.Wgt_2_781,.Wgt_2_782,.Wgt_2_783,.Wgt_2_784,
.Wgt_3_0,.Wgt_3_1,.Wgt_3_2,.Wgt_3_3,.Wgt_3_4,.Wgt_3_5,.Wgt_3_6,.Wgt_3_7,.Wgt_3_8,.Wgt_3_9,.Wgt_3_10,.Wgt_3_11,.Wgt_3_12,.Wgt_3_13,.Wgt_3_14,.Wgt_3_15,.Wgt_3_16,.Wgt_3_17,.Wgt_3_18,.Wgt_3_19,.Wgt_3_20,.Wgt_3_21,.Wgt_3_22,.Wgt_3_23,.Wgt_3_24,.Wgt_3_25,.Wgt_3_26,.Wgt_3_27,.Wgt_3_28,.Wgt_3_29,.Wgt_3_30,.Wgt_3_31,.Wgt_3_32,.Wgt_3_33,.Wgt_3_34,.Wgt_3_35,.Wgt_3_36,.Wgt_3_37,.Wgt_3_38,.Wgt_3_39,.Wgt_3_40,.Wgt_3_41,.Wgt_3_42,.Wgt_3_43,.Wgt_3_44,.Wgt_3_45,.Wgt_3_46,.Wgt_3_47,.Wgt_3_48,.Wgt_3_49,.Wgt_3_50,.Wgt_3_51,.Wgt_3_52,.Wgt_3_53,.Wgt_3_54,.Wgt_3_55,.Wgt_3_56,.Wgt_3_57,.Wgt_3_58,.Wgt_3_59,.Wgt_3_60,.Wgt_3_61,.Wgt_3_62,.Wgt_3_63,.Wgt_3_64,.Wgt_3_65,.Wgt_3_66,.Wgt_3_67,.Wgt_3_68,.Wgt_3_69,.Wgt_3_70,.Wgt_3_71,.Wgt_3_72,.Wgt_3_73,.Wgt_3_74,.Wgt_3_75,.Wgt_3_76,.Wgt_3_77,.Wgt_3_78,.Wgt_3_79,.Wgt_3_80,.Wgt_3_81,.Wgt_3_82,.Wgt_3_83,.Wgt_3_84,.Wgt_3_85,.Wgt_3_86,.Wgt_3_87,.Wgt_3_88,.Wgt_3_89,.Wgt_3_90,.Wgt_3_91,.Wgt_3_92,.Wgt_3_93,.Wgt_3_94,.Wgt_3_95,.Wgt_3_96,.Wgt_3_97,.Wgt_3_98,.Wgt_3_99,.Wgt_3_100,.Wgt_3_101,.Wgt_3_102,.Wgt_3_103,.Wgt_3_104,.Wgt_3_105,.Wgt_3_106,.Wgt_3_107,.Wgt_3_108,.Wgt_3_109,.Wgt_3_110,.Wgt_3_111,.Wgt_3_112,.Wgt_3_113,.Wgt_3_114,.Wgt_3_115,.Wgt_3_116,.Wgt_3_117,.Wgt_3_118,.Wgt_3_119,.Wgt_3_120,.Wgt_3_121,.Wgt_3_122,.Wgt_3_123,.Wgt_3_124,.Wgt_3_125,.Wgt_3_126,.Wgt_3_127,.Wgt_3_128,.Wgt_3_129,.Wgt_3_130,.Wgt_3_131,.Wgt_3_132,.Wgt_3_133,.Wgt_3_134,.Wgt_3_135,.Wgt_3_136,.Wgt_3_137,.Wgt_3_138,.Wgt_3_139,.Wgt_3_140,.Wgt_3_141,.Wgt_3_142,.Wgt_3_143,.Wgt_3_144,.Wgt_3_145,.Wgt_3_146,.Wgt_3_147,.Wgt_3_148,.Wgt_3_149,.Wgt_3_150,.Wgt_3_151,.Wgt_3_152,.Wgt_3_153,.Wgt_3_154,.Wgt_3_155,.Wgt_3_156,.Wgt_3_157,.Wgt_3_158,.Wgt_3_159,.Wgt_3_160,.Wgt_3_161,.Wgt_3_162,.Wgt_3_163,.Wgt_3_164,.Wgt_3_165,.Wgt_3_166,.Wgt_3_167,.Wgt_3_168,.Wgt_3_169,.Wgt_3_170,.Wgt_3_171,.Wgt_3_172,.Wgt_3_173,.Wgt_3_174,.Wgt_3_175,.Wgt_3_176,.Wgt_3_177,.Wgt_3_178,.Wgt_3_179,.Wgt_3_180,.Wgt_3_181,.Wgt_3_182,.Wgt_3_183,.Wgt_3_184,.Wgt_3_185,.Wgt_3_186,.Wgt_3_187,.Wgt_3_188,.Wgt_3_189,.Wgt_3_190,.Wgt_3_191,.Wgt_3_192,.Wgt_3_193,.Wgt_3_194,.Wgt_3_195,.Wgt_3_196,.Wgt_3_197,.Wgt_3_198,.Wgt_3_199,.Wgt_3_200,.Wgt_3_201,.Wgt_3_202,.Wgt_3_203,.Wgt_3_204,.Wgt_3_205,.Wgt_3_206,.Wgt_3_207,.Wgt_3_208,.Wgt_3_209,.Wgt_3_210,.Wgt_3_211,.Wgt_3_212,.Wgt_3_213,.Wgt_3_214,.Wgt_3_215,.Wgt_3_216,.Wgt_3_217,.Wgt_3_218,.Wgt_3_219,.Wgt_3_220,.Wgt_3_221,.Wgt_3_222,.Wgt_3_223,.Wgt_3_224,.Wgt_3_225,.Wgt_3_226,.Wgt_3_227,.Wgt_3_228,.Wgt_3_229,.Wgt_3_230,.Wgt_3_231,.Wgt_3_232,.Wgt_3_233,.Wgt_3_234,.Wgt_3_235,.Wgt_3_236,.Wgt_3_237,.Wgt_3_238,.Wgt_3_239,.Wgt_3_240,.Wgt_3_241,.Wgt_3_242,.Wgt_3_243,.Wgt_3_244,.Wgt_3_245,.Wgt_3_246,.Wgt_3_247,.Wgt_3_248,.Wgt_3_249,.Wgt_3_250,.Wgt_3_251,.Wgt_3_252,.Wgt_3_253,.Wgt_3_254,.Wgt_3_255,.Wgt_3_256,.Wgt_3_257,.Wgt_3_258,.Wgt_3_259,.Wgt_3_260,.Wgt_3_261,.Wgt_3_262,.Wgt_3_263,.Wgt_3_264,.Wgt_3_265,.Wgt_3_266,.Wgt_3_267,.Wgt_3_268,.Wgt_3_269,.Wgt_3_270,.Wgt_3_271,.Wgt_3_272,.Wgt_3_273,.Wgt_3_274,.Wgt_3_275,.Wgt_3_276,.Wgt_3_277,.Wgt_3_278,.Wgt_3_279,.Wgt_3_280,.Wgt_3_281,.Wgt_3_282,.Wgt_3_283,.Wgt_3_284,.Wgt_3_285,.Wgt_3_286,.Wgt_3_287,.Wgt_3_288,.Wgt_3_289,.Wgt_3_290,.Wgt_3_291,.Wgt_3_292,.Wgt_3_293,.Wgt_3_294,.Wgt_3_295,.Wgt_3_296,.Wgt_3_297,.Wgt_3_298,.Wgt_3_299,.Wgt_3_300,.Wgt_3_301,.Wgt_3_302,.Wgt_3_303,.Wgt_3_304,.Wgt_3_305,.Wgt_3_306,.Wgt_3_307,.Wgt_3_308,.Wgt_3_309,.Wgt_3_310,.Wgt_3_311,.Wgt_3_312,.Wgt_3_313,.Wgt_3_314,.Wgt_3_315,.Wgt_3_316,.Wgt_3_317,.Wgt_3_318,.Wgt_3_319,.Wgt_3_320,.Wgt_3_321,.Wgt_3_322,.Wgt_3_323,.Wgt_3_324,.Wgt_3_325,.Wgt_3_326,.Wgt_3_327,.Wgt_3_328,.Wgt_3_329,.Wgt_3_330,.Wgt_3_331,.Wgt_3_332,.Wgt_3_333,.Wgt_3_334,.Wgt_3_335,.Wgt_3_336,.Wgt_3_337,.Wgt_3_338,.Wgt_3_339,.Wgt_3_340,.Wgt_3_341,.Wgt_3_342,.Wgt_3_343,.Wgt_3_344,.Wgt_3_345,.Wgt_3_346,.Wgt_3_347,.Wgt_3_348,.Wgt_3_349,.Wgt_3_350,.Wgt_3_351,.Wgt_3_352,.Wgt_3_353,.Wgt_3_354,.Wgt_3_355,.Wgt_3_356,.Wgt_3_357,.Wgt_3_358,.Wgt_3_359,.Wgt_3_360,.Wgt_3_361,.Wgt_3_362,.Wgt_3_363,.Wgt_3_364,.Wgt_3_365,.Wgt_3_366,.Wgt_3_367,.Wgt_3_368,.Wgt_3_369,.Wgt_3_370,.Wgt_3_371,.Wgt_3_372,.Wgt_3_373,.Wgt_3_374,.Wgt_3_375,.Wgt_3_376,.Wgt_3_377,.Wgt_3_378,.Wgt_3_379,.Wgt_3_380,.Wgt_3_381,.Wgt_3_382,.Wgt_3_383,.Wgt_3_384,.Wgt_3_385,.Wgt_3_386,.Wgt_3_387,.Wgt_3_388,.Wgt_3_389,.Wgt_3_390,.Wgt_3_391,.Wgt_3_392,.Wgt_3_393,.Wgt_3_394,.Wgt_3_395,.Wgt_3_396,.Wgt_3_397,.Wgt_3_398,.Wgt_3_399,.Wgt_3_400,.Wgt_3_401,.Wgt_3_402,.Wgt_3_403,.Wgt_3_404,.Wgt_3_405,.Wgt_3_406,.Wgt_3_407,.Wgt_3_408,.Wgt_3_409,.Wgt_3_410,.Wgt_3_411,.Wgt_3_412,.Wgt_3_413,.Wgt_3_414,.Wgt_3_415,.Wgt_3_416,.Wgt_3_417,.Wgt_3_418,.Wgt_3_419,.Wgt_3_420,.Wgt_3_421,.Wgt_3_422,.Wgt_3_423,.Wgt_3_424,.Wgt_3_425,.Wgt_3_426,.Wgt_3_427,.Wgt_3_428,.Wgt_3_429,.Wgt_3_430,.Wgt_3_431,.Wgt_3_432,.Wgt_3_433,.Wgt_3_434,.Wgt_3_435,.Wgt_3_436,.Wgt_3_437,.Wgt_3_438,.Wgt_3_439,.Wgt_3_440,.Wgt_3_441,.Wgt_3_442,.Wgt_3_443,.Wgt_3_444,.Wgt_3_445,.Wgt_3_446,.Wgt_3_447,.Wgt_3_448,.Wgt_3_449,.Wgt_3_450,.Wgt_3_451,.Wgt_3_452,.Wgt_3_453,.Wgt_3_454,.Wgt_3_455,.Wgt_3_456,.Wgt_3_457,.Wgt_3_458,.Wgt_3_459,.Wgt_3_460,.Wgt_3_461,.Wgt_3_462,.Wgt_3_463,.Wgt_3_464,.Wgt_3_465,.Wgt_3_466,.Wgt_3_467,.Wgt_3_468,.Wgt_3_469,.Wgt_3_470,.Wgt_3_471,.Wgt_3_472,.Wgt_3_473,.Wgt_3_474,.Wgt_3_475,.Wgt_3_476,.Wgt_3_477,.Wgt_3_478,.Wgt_3_479,.Wgt_3_480,.Wgt_3_481,.Wgt_3_482,.Wgt_3_483,.Wgt_3_484,.Wgt_3_485,.Wgt_3_486,.Wgt_3_487,.Wgt_3_488,.Wgt_3_489,.Wgt_3_490,.Wgt_3_491,.Wgt_3_492,.Wgt_3_493,.Wgt_3_494,.Wgt_3_495,.Wgt_3_496,.Wgt_3_497,.Wgt_3_498,.Wgt_3_499,.Wgt_3_500,.Wgt_3_501,.Wgt_3_502,.Wgt_3_503,.Wgt_3_504,.Wgt_3_505,.Wgt_3_506,.Wgt_3_507,.Wgt_3_508,.Wgt_3_509,.Wgt_3_510,.Wgt_3_511,.Wgt_3_512,.Wgt_3_513,.Wgt_3_514,.Wgt_3_515,.Wgt_3_516,.Wgt_3_517,.Wgt_3_518,.Wgt_3_519,.Wgt_3_520,.Wgt_3_521,.Wgt_3_522,.Wgt_3_523,.Wgt_3_524,.Wgt_3_525,.Wgt_3_526,.Wgt_3_527,.Wgt_3_528,.Wgt_3_529,.Wgt_3_530,.Wgt_3_531,.Wgt_3_532,.Wgt_3_533,.Wgt_3_534,.Wgt_3_535,.Wgt_3_536,.Wgt_3_537,.Wgt_3_538,.Wgt_3_539,.Wgt_3_540,.Wgt_3_541,.Wgt_3_542,.Wgt_3_543,.Wgt_3_544,.Wgt_3_545,.Wgt_3_546,.Wgt_3_547,.Wgt_3_548,.Wgt_3_549,.Wgt_3_550,.Wgt_3_551,.Wgt_3_552,.Wgt_3_553,.Wgt_3_554,.Wgt_3_555,.Wgt_3_556,.Wgt_3_557,.Wgt_3_558,.Wgt_3_559,.Wgt_3_560,.Wgt_3_561,.Wgt_3_562,.Wgt_3_563,.Wgt_3_564,.Wgt_3_565,.Wgt_3_566,.Wgt_3_567,.Wgt_3_568,.Wgt_3_569,.Wgt_3_570,.Wgt_3_571,.Wgt_3_572,.Wgt_3_573,.Wgt_3_574,.Wgt_3_575,.Wgt_3_576,.Wgt_3_577,.Wgt_3_578,.Wgt_3_579,.Wgt_3_580,.Wgt_3_581,.Wgt_3_582,.Wgt_3_583,.Wgt_3_584,.Wgt_3_585,.Wgt_3_586,.Wgt_3_587,.Wgt_3_588,.Wgt_3_589,.Wgt_3_590,.Wgt_3_591,.Wgt_3_592,.Wgt_3_593,.Wgt_3_594,.Wgt_3_595,.Wgt_3_596,.Wgt_3_597,.Wgt_3_598,.Wgt_3_599,.Wgt_3_600,.Wgt_3_601,.Wgt_3_602,.Wgt_3_603,.Wgt_3_604,.Wgt_3_605,.Wgt_3_606,.Wgt_3_607,.Wgt_3_608,.Wgt_3_609,.Wgt_3_610,.Wgt_3_611,.Wgt_3_612,.Wgt_3_613,.Wgt_3_614,.Wgt_3_615,.Wgt_3_616,.Wgt_3_617,.Wgt_3_618,.Wgt_3_619,.Wgt_3_620,.Wgt_3_621,.Wgt_3_622,.Wgt_3_623,.Wgt_3_624,.Wgt_3_625,.Wgt_3_626,.Wgt_3_627,.Wgt_3_628,.Wgt_3_629,.Wgt_3_630,.Wgt_3_631,.Wgt_3_632,.Wgt_3_633,.Wgt_3_634,.Wgt_3_635,.Wgt_3_636,.Wgt_3_637,.Wgt_3_638,.Wgt_3_639,.Wgt_3_640,.Wgt_3_641,.Wgt_3_642,.Wgt_3_643,.Wgt_3_644,.Wgt_3_645,.Wgt_3_646,.Wgt_3_647,.Wgt_3_648,.Wgt_3_649,.Wgt_3_650,.Wgt_3_651,.Wgt_3_652,.Wgt_3_653,.Wgt_3_654,.Wgt_3_655,.Wgt_3_656,.Wgt_3_657,.Wgt_3_658,.Wgt_3_659,.Wgt_3_660,.Wgt_3_661,.Wgt_3_662,.Wgt_3_663,.Wgt_3_664,.Wgt_3_665,.Wgt_3_666,.Wgt_3_667,.Wgt_3_668,.Wgt_3_669,.Wgt_3_670,.Wgt_3_671,.Wgt_3_672,.Wgt_3_673,.Wgt_3_674,.Wgt_3_675,.Wgt_3_676,.Wgt_3_677,.Wgt_3_678,.Wgt_3_679,.Wgt_3_680,.Wgt_3_681,.Wgt_3_682,.Wgt_3_683,.Wgt_3_684,.Wgt_3_685,.Wgt_3_686,.Wgt_3_687,.Wgt_3_688,.Wgt_3_689,.Wgt_3_690,.Wgt_3_691,.Wgt_3_692,.Wgt_3_693,.Wgt_3_694,.Wgt_3_695,.Wgt_3_696,.Wgt_3_697,.Wgt_3_698,.Wgt_3_699,.Wgt_3_700,.Wgt_3_701,.Wgt_3_702,.Wgt_3_703,.Wgt_3_704,.Wgt_3_705,.Wgt_3_706,.Wgt_3_707,.Wgt_3_708,.Wgt_3_709,.Wgt_3_710,.Wgt_3_711,.Wgt_3_712,.Wgt_3_713,.Wgt_3_714,.Wgt_3_715,.Wgt_3_716,.Wgt_3_717,.Wgt_3_718,.Wgt_3_719,.Wgt_3_720,.Wgt_3_721,.Wgt_3_722,.Wgt_3_723,.Wgt_3_724,.Wgt_3_725,.Wgt_3_726,.Wgt_3_727,.Wgt_3_728,.Wgt_3_729,.Wgt_3_730,.Wgt_3_731,.Wgt_3_732,.Wgt_3_733,.Wgt_3_734,.Wgt_3_735,.Wgt_3_736,.Wgt_3_737,.Wgt_3_738,.Wgt_3_739,.Wgt_3_740,.Wgt_3_741,.Wgt_3_742,.Wgt_3_743,.Wgt_3_744,.Wgt_3_745,.Wgt_3_746,.Wgt_3_747,.Wgt_3_748,.Wgt_3_749,.Wgt_3_750,.Wgt_3_751,.Wgt_3_752,.Wgt_3_753,.Wgt_3_754,.Wgt_3_755,.Wgt_3_756,.Wgt_3_757,.Wgt_3_758,.Wgt_3_759,.Wgt_3_760,.Wgt_3_761,.Wgt_3_762,.Wgt_3_763,.Wgt_3_764,.Wgt_3_765,.Wgt_3_766,.Wgt_3_767,.Wgt_3_768,.Wgt_3_769,.Wgt_3_770,.Wgt_3_771,.Wgt_3_772,.Wgt_3_773,.Wgt_3_774,.Wgt_3_775,.Wgt_3_776,.Wgt_3_777,.Wgt_3_778,.Wgt_3_779,.Wgt_3_780,.Wgt_3_781,.Wgt_3_782,.Wgt_3_783,.Wgt_3_784,
.Wgt_4_0,.Wgt_4_1,.Wgt_4_2,.Wgt_4_3,.Wgt_4_4,.Wgt_4_5,.Wgt_4_6,.Wgt_4_7,.Wgt_4_8,.Wgt_4_9,.Wgt_4_10,.Wgt_4_11,.Wgt_4_12,.Wgt_4_13,.Wgt_4_14,.Wgt_4_15,.Wgt_4_16,.Wgt_4_17,.Wgt_4_18,.Wgt_4_19,.Wgt_4_20,.Wgt_4_21,.Wgt_4_22,.Wgt_4_23,.Wgt_4_24,.Wgt_4_25,.Wgt_4_26,.Wgt_4_27,.Wgt_4_28,.Wgt_4_29,.Wgt_4_30,.Wgt_4_31,.Wgt_4_32,.Wgt_4_33,.Wgt_4_34,.Wgt_4_35,.Wgt_4_36,.Wgt_4_37,.Wgt_4_38,.Wgt_4_39,.Wgt_4_40,.Wgt_4_41,.Wgt_4_42,.Wgt_4_43,.Wgt_4_44,.Wgt_4_45,.Wgt_4_46,.Wgt_4_47,.Wgt_4_48,.Wgt_4_49,.Wgt_4_50,.Wgt_4_51,.Wgt_4_52,.Wgt_4_53,.Wgt_4_54,.Wgt_4_55,.Wgt_4_56,.Wgt_4_57,.Wgt_4_58,.Wgt_4_59,.Wgt_4_60,.Wgt_4_61,.Wgt_4_62,.Wgt_4_63,.Wgt_4_64,.Wgt_4_65,.Wgt_4_66,.Wgt_4_67,.Wgt_4_68,.Wgt_4_69,.Wgt_4_70,.Wgt_4_71,.Wgt_4_72,.Wgt_4_73,.Wgt_4_74,.Wgt_4_75,.Wgt_4_76,.Wgt_4_77,.Wgt_4_78,.Wgt_4_79,.Wgt_4_80,.Wgt_4_81,.Wgt_4_82,.Wgt_4_83,.Wgt_4_84,.Wgt_4_85,.Wgt_4_86,.Wgt_4_87,.Wgt_4_88,.Wgt_4_89,.Wgt_4_90,.Wgt_4_91,.Wgt_4_92,.Wgt_4_93,.Wgt_4_94,.Wgt_4_95,.Wgt_4_96,.Wgt_4_97,.Wgt_4_98,.Wgt_4_99,.Wgt_4_100,.Wgt_4_101,.Wgt_4_102,.Wgt_4_103,.Wgt_4_104,.Wgt_4_105,.Wgt_4_106,.Wgt_4_107,.Wgt_4_108,.Wgt_4_109,.Wgt_4_110,.Wgt_4_111,.Wgt_4_112,.Wgt_4_113,.Wgt_4_114,.Wgt_4_115,.Wgt_4_116,.Wgt_4_117,.Wgt_4_118,.Wgt_4_119,.Wgt_4_120,.Wgt_4_121,.Wgt_4_122,.Wgt_4_123,.Wgt_4_124,.Wgt_4_125,.Wgt_4_126,.Wgt_4_127,.Wgt_4_128,.Wgt_4_129,.Wgt_4_130,.Wgt_4_131,.Wgt_4_132,.Wgt_4_133,.Wgt_4_134,.Wgt_4_135,.Wgt_4_136,.Wgt_4_137,.Wgt_4_138,.Wgt_4_139,.Wgt_4_140,.Wgt_4_141,.Wgt_4_142,.Wgt_4_143,.Wgt_4_144,.Wgt_4_145,.Wgt_4_146,.Wgt_4_147,.Wgt_4_148,.Wgt_4_149,.Wgt_4_150,.Wgt_4_151,.Wgt_4_152,.Wgt_4_153,.Wgt_4_154,.Wgt_4_155,.Wgt_4_156,.Wgt_4_157,.Wgt_4_158,.Wgt_4_159,.Wgt_4_160,.Wgt_4_161,.Wgt_4_162,.Wgt_4_163,.Wgt_4_164,.Wgt_4_165,.Wgt_4_166,.Wgt_4_167,.Wgt_4_168,.Wgt_4_169,.Wgt_4_170,.Wgt_4_171,.Wgt_4_172,.Wgt_4_173,.Wgt_4_174,.Wgt_4_175,.Wgt_4_176,.Wgt_4_177,.Wgt_4_178,.Wgt_4_179,.Wgt_4_180,.Wgt_4_181,.Wgt_4_182,.Wgt_4_183,.Wgt_4_184,.Wgt_4_185,.Wgt_4_186,.Wgt_4_187,.Wgt_4_188,.Wgt_4_189,.Wgt_4_190,.Wgt_4_191,.Wgt_4_192,.Wgt_4_193,.Wgt_4_194,.Wgt_4_195,.Wgt_4_196,.Wgt_4_197,.Wgt_4_198,.Wgt_4_199,.Wgt_4_200,.Wgt_4_201,.Wgt_4_202,.Wgt_4_203,.Wgt_4_204,.Wgt_4_205,.Wgt_4_206,.Wgt_4_207,.Wgt_4_208,.Wgt_4_209,.Wgt_4_210,.Wgt_4_211,.Wgt_4_212,.Wgt_4_213,.Wgt_4_214,.Wgt_4_215,.Wgt_4_216,.Wgt_4_217,.Wgt_4_218,.Wgt_4_219,.Wgt_4_220,.Wgt_4_221,.Wgt_4_222,.Wgt_4_223,.Wgt_4_224,.Wgt_4_225,.Wgt_4_226,.Wgt_4_227,.Wgt_4_228,.Wgt_4_229,.Wgt_4_230,.Wgt_4_231,.Wgt_4_232,.Wgt_4_233,.Wgt_4_234,.Wgt_4_235,.Wgt_4_236,.Wgt_4_237,.Wgt_4_238,.Wgt_4_239,.Wgt_4_240,.Wgt_4_241,.Wgt_4_242,.Wgt_4_243,.Wgt_4_244,.Wgt_4_245,.Wgt_4_246,.Wgt_4_247,.Wgt_4_248,.Wgt_4_249,.Wgt_4_250,.Wgt_4_251,.Wgt_4_252,.Wgt_4_253,.Wgt_4_254,.Wgt_4_255,.Wgt_4_256,.Wgt_4_257,.Wgt_4_258,.Wgt_4_259,.Wgt_4_260,.Wgt_4_261,.Wgt_4_262,.Wgt_4_263,.Wgt_4_264,.Wgt_4_265,.Wgt_4_266,.Wgt_4_267,.Wgt_4_268,.Wgt_4_269,.Wgt_4_270,.Wgt_4_271,.Wgt_4_272,.Wgt_4_273,.Wgt_4_274,.Wgt_4_275,.Wgt_4_276,.Wgt_4_277,.Wgt_4_278,.Wgt_4_279,.Wgt_4_280,.Wgt_4_281,.Wgt_4_282,.Wgt_4_283,.Wgt_4_284,.Wgt_4_285,.Wgt_4_286,.Wgt_4_287,.Wgt_4_288,.Wgt_4_289,.Wgt_4_290,.Wgt_4_291,.Wgt_4_292,.Wgt_4_293,.Wgt_4_294,.Wgt_4_295,.Wgt_4_296,.Wgt_4_297,.Wgt_4_298,.Wgt_4_299,.Wgt_4_300,.Wgt_4_301,.Wgt_4_302,.Wgt_4_303,.Wgt_4_304,.Wgt_4_305,.Wgt_4_306,.Wgt_4_307,.Wgt_4_308,.Wgt_4_309,.Wgt_4_310,.Wgt_4_311,.Wgt_4_312,.Wgt_4_313,.Wgt_4_314,.Wgt_4_315,.Wgt_4_316,.Wgt_4_317,.Wgt_4_318,.Wgt_4_319,.Wgt_4_320,.Wgt_4_321,.Wgt_4_322,.Wgt_4_323,.Wgt_4_324,.Wgt_4_325,.Wgt_4_326,.Wgt_4_327,.Wgt_4_328,.Wgt_4_329,.Wgt_4_330,.Wgt_4_331,.Wgt_4_332,.Wgt_4_333,.Wgt_4_334,.Wgt_4_335,.Wgt_4_336,.Wgt_4_337,.Wgt_4_338,.Wgt_4_339,.Wgt_4_340,.Wgt_4_341,.Wgt_4_342,.Wgt_4_343,.Wgt_4_344,.Wgt_4_345,.Wgt_4_346,.Wgt_4_347,.Wgt_4_348,.Wgt_4_349,.Wgt_4_350,.Wgt_4_351,.Wgt_4_352,.Wgt_4_353,.Wgt_4_354,.Wgt_4_355,.Wgt_4_356,.Wgt_4_357,.Wgt_4_358,.Wgt_4_359,.Wgt_4_360,.Wgt_4_361,.Wgt_4_362,.Wgt_4_363,.Wgt_4_364,.Wgt_4_365,.Wgt_4_366,.Wgt_4_367,.Wgt_4_368,.Wgt_4_369,.Wgt_4_370,.Wgt_4_371,.Wgt_4_372,.Wgt_4_373,.Wgt_4_374,.Wgt_4_375,.Wgt_4_376,.Wgt_4_377,.Wgt_4_378,.Wgt_4_379,.Wgt_4_380,.Wgt_4_381,.Wgt_4_382,.Wgt_4_383,.Wgt_4_384,.Wgt_4_385,.Wgt_4_386,.Wgt_4_387,.Wgt_4_388,.Wgt_4_389,.Wgt_4_390,.Wgt_4_391,.Wgt_4_392,.Wgt_4_393,.Wgt_4_394,.Wgt_4_395,.Wgt_4_396,.Wgt_4_397,.Wgt_4_398,.Wgt_4_399,.Wgt_4_400,.Wgt_4_401,.Wgt_4_402,.Wgt_4_403,.Wgt_4_404,.Wgt_4_405,.Wgt_4_406,.Wgt_4_407,.Wgt_4_408,.Wgt_4_409,.Wgt_4_410,.Wgt_4_411,.Wgt_4_412,.Wgt_4_413,.Wgt_4_414,.Wgt_4_415,.Wgt_4_416,.Wgt_4_417,.Wgt_4_418,.Wgt_4_419,.Wgt_4_420,.Wgt_4_421,.Wgt_4_422,.Wgt_4_423,.Wgt_4_424,.Wgt_4_425,.Wgt_4_426,.Wgt_4_427,.Wgt_4_428,.Wgt_4_429,.Wgt_4_430,.Wgt_4_431,.Wgt_4_432,.Wgt_4_433,.Wgt_4_434,.Wgt_4_435,.Wgt_4_436,.Wgt_4_437,.Wgt_4_438,.Wgt_4_439,.Wgt_4_440,.Wgt_4_441,.Wgt_4_442,.Wgt_4_443,.Wgt_4_444,.Wgt_4_445,.Wgt_4_446,.Wgt_4_447,.Wgt_4_448,.Wgt_4_449,.Wgt_4_450,.Wgt_4_451,.Wgt_4_452,.Wgt_4_453,.Wgt_4_454,.Wgt_4_455,.Wgt_4_456,.Wgt_4_457,.Wgt_4_458,.Wgt_4_459,.Wgt_4_460,.Wgt_4_461,.Wgt_4_462,.Wgt_4_463,.Wgt_4_464,.Wgt_4_465,.Wgt_4_466,.Wgt_4_467,.Wgt_4_468,.Wgt_4_469,.Wgt_4_470,.Wgt_4_471,.Wgt_4_472,.Wgt_4_473,.Wgt_4_474,.Wgt_4_475,.Wgt_4_476,.Wgt_4_477,.Wgt_4_478,.Wgt_4_479,.Wgt_4_480,.Wgt_4_481,.Wgt_4_482,.Wgt_4_483,.Wgt_4_484,.Wgt_4_485,.Wgt_4_486,.Wgt_4_487,.Wgt_4_488,.Wgt_4_489,.Wgt_4_490,.Wgt_4_491,.Wgt_4_492,.Wgt_4_493,.Wgt_4_494,.Wgt_4_495,.Wgt_4_496,.Wgt_4_497,.Wgt_4_498,.Wgt_4_499,.Wgt_4_500,.Wgt_4_501,.Wgt_4_502,.Wgt_4_503,.Wgt_4_504,.Wgt_4_505,.Wgt_4_506,.Wgt_4_507,.Wgt_4_508,.Wgt_4_509,.Wgt_4_510,.Wgt_4_511,.Wgt_4_512,.Wgt_4_513,.Wgt_4_514,.Wgt_4_515,.Wgt_4_516,.Wgt_4_517,.Wgt_4_518,.Wgt_4_519,.Wgt_4_520,.Wgt_4_521,.Wgt_4_522,.Wgt_4_523,.Wgt_4_524,.Wgt_4_525,.Wgt_4_526,.Wgt_4_527,.Wgt_4_528,.Wgt_4_529,.Wgt_4_530,.Wgt_4_531,.Wgt_4_532,.Wgt_4_533,.Wgt_4_534,.Wgt_4_535,.Wgt_4_536,.Wgt_4_537,.Wgt_4_538,.Wgt_4_539,.Wgt_4_540,.Wgt_4_541,.Wgt_4_542,.Wgt_4_543,.Wgt_4_544,.Wgt_4_545,.Wgt_4_546,.Wgt_4_547,.Wgt_4_548,.Wgt_4_549,.Wgt_4_550,.Wgt_4_551,.Wgt_4_552,.Wgt_4_553,.Wgt_4_554,.Wgt_4_555,.Wgt_4_556,.Wgt_4_557,.Wgt_4_558,.Wgt_4_559,.Wgt_4_560,.Wgt_4_561,.Wgt_4_562,.Wgt_4_563,.Wgt_4_564,.Wgt_4_565,.Wgt_4_566,.Wgt_4_567,.Wgt_4_568,.Wgt_4_569,.Wgt_4_570,.Wgt_4_571,.Wgt_4_572,.Wgt_4_573,.Wgt_4_574,.Wgt_4_575,.Wgt_4_576,.Wgt_4_577,.Wgt_4_578,.Wgt_4_579,.Wgt_4_580,.Wgt_4_581,.Wgt_4_582,.Wgt_4_583,.Wgt_4_584,.Wgt_4_585,.Wgt_4_586,.Wgt_4_587,.Wgt_4_588,.Wgt_4_589,.Wgt_4_590,.Wgt_4_591,.Wgt_4_592,.Wgt_4_593,.Wgt_4_594,.Wgt_4_595,.Wgt_4_596,.Wgt_4_597,.Wgt_4_598,.Wgt_4_599,.Wgt_4_600,.Wgt_4_601,.Wgt_4_602,.Wgt_4_603,.Wgt_4_604,.Wgt_4_605,.Wgt_4_606,.Wgt_4_607,.Wgt_4_608,.Wgt_4_609,.Wgt_4_610,.Wgt_4_611,.Wgt_4_612,.Wgt_4_613,.Wgt_4_614,.Wgt_4_615,.Wgt_4_616,.Wgt_4_617,.Wgt_4_618,.Wgt_4_619,.Wgt_4_620,.Wgt_4_621,.Wgt_4_622,.Wgt_4_623,.Wgt_4_624,.Wgt_4_625,.Wgt_4_626,.Wgt_4_627,.Wgt_4_628,.Wgt_4_629,.Wgt_4_630,.Wgt_4_631,.Wgt_4_632,.Wgt_4_633,.Wgt_4_634,.Wgt_4_635,.Wgt_4_636,.Wgt_4_637,.Wgt_4_638,.Wgt_4_639,.Wgt_4_640,.Wgt_4_641,.Wgt_4_642,.Wgt_4_643,.Wgt_4_644,.Wgt_4_645,.Wgt_4_646,.Wgt_4_647,.Wgt_4_648,.Wgt_4_649,.Wgt_4_650,.Wgt_4_651,.Wgt_4_652,.Wgt_4_653,.Wgt_4_654,.Wgt_4_655,.Wgt_4_656,.Wgt_4_657,.Wgt_4_658,.Wgt_4_659,.Wgt_4_660,.Wgt_4_661,.Wgt_4_662,.Wgt_4_663,.Wgt_4_664,.Wgt_4_665,.Wgt_4_666,.Wgt_4_667,.Wgt_4_668,.Wgt_4_669,.Wgt_4_670,.Wgt_4_671,.Wgt_4_672,.Wgt_4_673,.Wgt_4_674,.Wgt_4_675,.Wgt_4_676,.Wgt_4_677,.Wgt_4_678,.Wgt_4_679,.Wgt_4_680,.Wgt_4_681,.Wgt_4_682,.Wgt_4_683,.Wgt_4_684,.Wgt_4_685,.Wgt_4_686,.Wgt_4_687,.Wgt_4_688,.Wgt_4_689,.Wgt_4_690,.Wgt_4_691,.Wgt_4_692,.Wgt_4_693,.Wgt_4_694,.Wgt_4_695,.Wgt_4_696,.Wgt_4_697,.Wgt_4_698,.Wgt_4_699,.Wgt_4_700,.Wgt_4_701,.Wgt_4_702,.Wgt_4_703,.Wgt_4_704,.Wgt_4_705,.Wgt_4_706,.Wgt_4_707,.Wgt_4_708,.Wgt_4_709,.Wgt_4_710,.Wgt_4_711,.Wgt_4_712,.Wgt_4_713,.Wgt_4_714,.Wgt_4_715,.Wgt_4_716,.Wgt_4_717,.Wgt_4_718,.Wgt_4_719,.Wgt_4_720,.Wgt_4_721,.Wgt_4_722,.Wgt_4_723,.Wgt_4_724,.Wgt_4_725,.Wgt_4_726,.Wgt_4_727,.Wgt_4_728,.Wgt_4_729,.Wgt_4_730,.Wgt_4_731,.Wgt_4_732,.Wgt_4_733,.Wgt_4_734,.Wgt_4_735,.Wgt_4_736,.Wgt_4_737,.Wgt_4_738,.Wgt_4_739,.Wgt_4_740,.Wgt_4_741,.Wgt_4_742,.Wgt_4_743,.Wgt_4_744,.Wgt_4_745,.Wgt_4_746,.Wgt_4_747,.Wgt_4_748,.Wgt_4_749,.Wgt_4_750,.Wgt_4_751,.Wgt_4_752,.Wgt_4_753,.Wgt_4_754,.Wgt_4_755,.Wgt_4_756,.Wgt_4_757,.Wgt_4_758,.Wgt_4_759,.Wgt_4_760,.Wgt_4_761,.Wgt_4_762,.Wgt_4_763,.Wgt_4_764,.Wgt_4_765,.Wgt_4_766,.Wgt_4_767,.Wgt_4_768,.Wgt_4_769,.Wgt_4_770,.Wgt_4_771,.Wgt_4_772,.Wgt_4_773,.Wgt_4_774,.Wgt_4_775,.Wgt_4_776,.Wgt_4_777,.Wgt_4_778,.Wgt_4_779,.Wgt_4_780,.Wgt_4_781,.Wgt_4_782,.Wgt_4_783,.Wgt_4_784,
.Wgt_5_0,.Wgt_5_1,.Wgt_5_2,.Wgt_5_3,.Wgt_5_4,.Wgt_5_5,.Wgt_5_6,.Wgt_5_7,.Wgt_5_8,.Wgt_5_9,.Wgt_5_10,.Wgt_5_11,.Wgt_5_12,.Wgt_5_13,.Wgt_5_14,.Wgt_5_15,.Wgt_5_16,.Wgt_5_17,.Wgt_5_18,.Wgt_5_19,.Wgt_5_20,.Wgt_5_21,.Wgt_5_22,.Wgt_5_23,.Wgt_5_24,.Wgt_5_25,.Wgt_5_26,.Wgt_5_27,.Wgt_5_28,.Wgt_5_29,.Wgt_5_30,.Wgt_5_31,.Wgt_5_32,.Wgt_5_33,.Wgt_5_34,.Wgt_5_35,.Wgt_5_36,.Wgt_5_37,.Wgt_5_38,.Wgt_5_39,.Wgt_5_40,.Wgt_5_41,.Wgt_5_42,.Wgt_5_43,.Wgt_5_44,.Wgt_5_45,.Wgt_5_46,.Wgt_5_47,.Wgt_5_48,.Wgt_5_49,.Wgt_5_50,.Wgt_5_51,.Wgt_5_52,.Wgt_5_53,.Wgt_5_54,.Wgt_5_55,.Wgt_5_56,.Wgt_5_57,.Wgt_5_58,.Wgt_5_59,.Wgt_5_60,.Wgt_5_61,.Wgt_5_62,.Wgt_5_63,.Wgt_5_64,.Wgt_5_65,.Wgt_5_66,.Wgt_5_67,.Wgt_5_68,.Wgt_5_69,.Wgt_5_70,.Wgt_5_71,.Wgt_5_72,.Wgt_5_73,.Wgt_5_74,.Wgt_5_75,.Wgt_5_76,.Wgt_5_77,.Wgt_5_78,.Wgt_5_79,.Wgt_5_80,.Wgt_5_81,.Wgt_5_82,.Wgt_5_83,.Wgt_5_84,.Wgt_5_85,.Wgt_5_86,.Wgt_5_87,.Wgt_5_88,.Wgt_5_89,.Wgt_5_90,.Wgt_5_91,.Wgt_5_92,.Wgt_5_93,.Wgt_5_94,.Wgt_5_95,.Wgt_5_96,.Wgt_5_97,.Wgt_5_98,.Wgt_5_99,.Wgt_5_100,.Wgt_5_101,.Wgt_5_102,.Wgt_5_103,.Wgt_5_104,.Wgt_5_105,.Wgt_5_106,.Wgt_5_107,.Wgt_5_108,.Wgt_5_109,.Wgt_5_110,.Wgt_5_111,.Wgt_5_112,.Wgt_5_113,.Wgt_5_114,.Wgt_5_115,.Wgt_5_116,.Wgt_5_117,.Wgt_5_118,.Wgt_5_119,.Wgt_5_120,.Wgt_5_121,.Wgt_5_122,.Wgt_5_123,.Wgt_5_124,.Wgt_5_125,.Wgt_5_126,.Wgt_5_127,.Wgt_5_128,.Wgt_5_129,.Wgt_5_130,.Wgt_5_131,.Wgt_5_132,.Wgt_5_133,.Wgt_5_134,.Wgt_5_135,.Wgt_5_136,.Wgt_5_137,.Wgt_5_138,.Wgt_5_139,.Wgt_5_140,.Wgt_5_141,.Wgt_5_142,.Wgt_5_143,.Wgt_5_144,.Wgt_5_145,.Wgt_5_146,.Wgt_5_147,.Wgt_5_148,.Wgt_5_149,.Wgt_5_150,.Wgt_5_151,.Wgt_5_152,.Wgt_5_153,.Wgt_5_154,.Wgt_5_155,.Wgt_5_156,.Wgt_5_157,.Wgt_5_158,.Wgt_5_159,.Wgt_5_160,.Wgt_5_161,.Wgt_5_162,.Wgt_5_163,.Wgt_5_164,.Wgt_5_165,.Wgt_5_166,.Wgt_5_167,.Wgt_5_168,.Wgt_5_169,.Wgt_5_170,.Wgt_5_171,.Wgt_5_172,.Wgt_5_173,.Wgt_5_174,.Wgt_5_175,.Wgt_5_176,.Wgt_5_177,.Wgt_5_178,.Wgt_5_179,.Wgt_5_180,.Wgt_5_181,.Wgt_5_182,.Wgt_5_183,.Wgt_5_184,.Wgt_5_185,.Wgt_5_186,.Wgt_5_187,.Wgt_5_188,.Wgt_5_189,.Wgt_5_190,.Wgt_5_191,.Wgt_5_192,.Wgt_5_193,.Wgt_5_194,.Wgt_5_195,.Wgt_5_196,.Wgt_5_197,.Wgt_5_198,.Wgt_5_199,.Wgt_5_200,.Wgt_5_201,.Wgt_5_202,.Wgt_5_203,.Wgt_5_204,.Wgt_5_205,.Wgt_5_206,.Wgt_5_207,.Wgt_5_208,.Wgt_5_209,.Wgt_5_210,.Wgt_5_211,.Wgt_5_212,.Wgt_5_213,.Wgt_5_214,.Wgt_5_215,.Wgt_5_216,.Wgt_5_217,.Wgt_5_218,.Wgt_5_219,.Wgt_5_220,.Wgt_5_221,.Wgt_5_222,.Wgt_5_223,.Wgt_5_224,.Wgt_5_225,.Wgt_5_226,.Wgt_5_227,.Wgt_5_228,.Wgt_5_229,.Wgt_5_230,.Wgt_5_231,.Wgt_5_232,.Wgt_5_233,.Wgt_5_234,.Wgt_5_235,.Wgt_5_236,.Wgt_5_237,.Wgt_5_238,.Wgt_5_239,.Wgt_5_240,.Wgt_5_241,.Wgt_5_242,.Wgt_5_243,.Wgt_5_244,.Wgt_5_245,.Wgt_5_246,.Wgt_5_247,.Wgt_5_248,.Wgt_5_249,.Wgt_5_250,.Wgt_5_251,.Wgt_5_252,.Wgt_5_253,.Wgt_5_254,.Wgt_5_255,.Wgt_5_256,.Wgt_5_257,.Wgt_5_258,.Wgt_5_259,.Wgt_5_260,.Wgt_5_261,.Wgt_5_262,.Wgt_5_263,.Wgt_5_264,.Wgt_5_265,.Wgt_5_266,.Wgt_5_267,.Wgt_5_268,.Wgt_5_269,.Wgt_5_270,.Wgt_5_271,.Wgt_5_272,.Wgt_5_273,.Wgt_5_274,.Wgt_5_275,.Wgt_5_276,.Wgt_5_277,.Wgt_5_278,.Wgt_5_279,.Wgt_5_280,.Wgt_5_281,.Wgt_5_282,.Wgt_5_283,.Wgt_5_284,.Wgt_5_285,.Wgt_5_286,.Wgt_5_287,.Wgt_5_288,.Wgt_5_289,.Wgt_5_290,.Wgt_5_291,.Wgt_5_292,.Wgt_5_293,.Wgt_5_294,.Wgt_5_295,.Wgt_5_296,.Wgt_5_297,.Wgt_5_298,.Wgt_5_299,.Wgt_5_300,.Wgt_5_301,.Wgt_5_302,.Wgt_5_303,.Wgt_5_304,.Wgt_5_305,.Wgt_5_306,.Wgt_5_307,.Wgt_5_308,.Wgt_5_309,.Wgt_5_310,.Wgt_5_311,.Wgt_5_312,.Wgt_5_313,.Wgt_5_314,.Wgt_5_315,.Wgt_5_316,.Wgt_5_317,.Wgt_5_318,.Wgt_5_319,.Wgt_5_320,.Wgt_5_321,.Wgt_5_322,.Wgt_5_323,.Wgt_5_324,.Wgt_5_325,.Wgt_5_326,.Wgt_5_327,.Wgt_5_328,.Wgt_5_329,.Wgt_5_330,.Wgt_5_331,.Wgt_5_332,.Wgt_5_333,.Wgt_5_334,.Wgt_5_335,.Wgt_5_336,.Wgt_5_337,.Wgt_5_338,.Wgt_5_339,.Wgt_5_340,.Wgt_5_341,.Wgt_5_342,.Wgt_5_343,.Wgt_5_344,.Wgt_5_345,.Wgt_5_346,.Wgt_5_347,.Wgt_5_348,.Wgt_5_349,.Wgt_5_350,.Wgt_5_351,.Wgt_5_352,.Wgt_5_353,.Wgt_5_354,.Wgt_5_355,.Wgt_5_356,.Wgt_5_357,.Wgt_5_358,.Wgt_5_359,.Wgt_5_360,.Wgt_5_361,.Wgt_5_362,.Wgt_5_363,.Wgt_5_364,.Wgt_5_365,.Wgt_5_366,.Wgt_5_367,.Wgt_5_368,.Wgt_5_369,.Wgt_5_370,.Wgt_5_371,.Wgt_5_372,.Wgt_5_373,.Wgt_5_374,.Wgt_5_375,.Wgt_5_376,.Wgt_5_377,.Wgt_5_378,.Wgt_5_379,.Wgt_5_380,.Wgt_5_381,.Wgt_5_382,.Wgt_5_383,.Wgt_5_384,.Wgt_5_385,.Wgt_5_386,.Wgt_5_387,.Wgt_5_388,.Wgt_5_389,.Wgt_5_390,.Wgt_5_391,.Wgt_5_392,.Wgt_5_393,.Wgt_5_394,.Wgt_5_395,.Wgt_5_396,.Wgt_5_397,.Wgt_5_398,.Wgt_5_399,.Wgt_5_400,.Wgt_5_401,.Wgt_5_402,.Wgt_5_403,.Wgt_5_404,.Wgt_5_405,.Wgt_5_406,.Wgt_5_407,.Wgt_5_408,.Wgt_5_409,.Wgt_5_410,.Wgt_5_411,.Wgt_5_412,.Wgt_5_413,.Wgt_5_414,.Wgt_5_415,.Wgt_5_416,.Wgt_5_417,.Wgt_5_418,.Wgt_5_419,.Wgt_5_420,.Wgt_5_421,.Wgt_5_422,.Wgt_5_423,.Wgt_5_424,.Wgt_5_425,.Wgt_5_426,.Wgt_5_427,.Wgt_5_428,.Wgt_5_429,.Wgt_5_430,.Wgt_5_431,.Wgt_5_432,.Wgt_5_433,.Wgt_5_434,.Wgt_5_435,.Wgt_5_436,.Wgt_5_437,.Wgt_5_438,.Wgt_5_439,.Wgt_5_440,.Wgt_5_441,.Wgt_5_442,.Wgt_5_443,.Wgt_5_444,.Wgt_5_445,.Wgt_5_446,.Wgt_5_447,.Wgt_5_448,.Wgt_5_449,.Wgt_5_450,.Wgt_5_451,.Wgt_5_452,.Wgt_5_453,.Wgt_5_454,.Wgt_5_455,.Wgt_5_456,.Wgt_5_457,.Wgt_5_458,.Wgt_5_459,.Wgt_5_460,.Wgt_5_461,.Wgt_5_462,.Wgt_5_463,.Wgt_5_464,.Wgt_5_465,.Wgt_5_466,.Wgt_5_467,.Wgt_5_468,.Wgt_5_469,.Wgt_5_470,.Wgt_5_471,.Wgt_5_472,.Wgt_5_473,.Wgt_5_474,.Wgt_5_475,.Wgt_5_476,.Wgt_5_477,.Wgt_5_478,.Wgt_5_479,.Wgt_5_480,.Wgt_5_481,.Wgt_5_482,.Wgt_5_483,.Wgt_5_484,.Wgt_5_485,.Wgt_5_486,.Wgt_5_487,.Wgt_5_488,.Wgt_5_489,.Wgt_5_490,.Wgt_5_491,.Wgt_5_492,.Wgt_5_493,.Wgt_5_494,.Wgt_5_495,.Wgt_5_496,.Wgt_5_497,.Wgt_5_498,.Wgt_5_499,.Wgt_5_500,.Wgt_5_501,.Wgt_5_502,.Wgt_5_503,.Wgt_5_504,.Wgt_5_505,.Wgt_5_506,.Wgt_5_507,.Wgt_5_508,.Wgt_5_509,.Wgt_5_510,.Wgt_5_511,.Wgt_5_512,.Wgt_5_513,.Wgt_5_514,.Wgt_5_515,.Wgt_5_516,.Wgt_5_517,.Wgt_5_518,.Wgt_5_519,.Wgt_5_520,.Wgt_5_521,.Wgt_5_522,.Wgt_5_523,.Wgt_5_524,.Wgt_5_525,.Wgt_5_526,.Wgt_5_527,.Wgt_5_528,.Wgt_5_529,.Wgt_5_530,.Wgt_5_531,.Wgt_5_532,.Wgt_5_533,.Wgt_5_534,.Wgt_5_535,.Wgt_5_536,.Wgt_5_537,.Wgt_5_538,.Wgt_5_539,.Wgt_5_540,.Wgt_5_541,.Wgt_5_542,.Wgt_5_543,.Wgt_5_544,.Wgt_5_545,.Wgt_5_546,.Wgt_5_547,.Wgt_5_548,.Wgt_5_549,.Wgt_5_550,.Wgt_5_551,.Wgt_5_552,.Wgt_5_553,.Wgt_5_554,.Wgt_5_555,.Wgt_5_556,.Wgt_5_557,.Wgt_5_558,.Wgt_5_559,.Wgt_5_560,.Wgt_5_561,.Wgt_5_562,.Wgt_5_563,.Wgt_5_564,.Wgt_5_565,.Wgt_5_566,.Wgt_5_567,.Wgt_5_568,.Wgt_5_569,.Wgt_5_570,.Wgt_5_571,.Wgt_5_572,.Wgt_5_573,.Wgt_5_574,.Wgt_5_575,.Wgt_5_576,.Wgt_5_577,.Wgt_5_578,.Wgt_5_579,.Wgt_5_580,.Wgt_5_581,.Wgt_5_582,.Wgt_5_583,.Wgt_5_584,.Wgt_5_585,.Wgt_5_586,.Wgt_5_587,.Wgt_5_588,.Wgt_5_589,.Wgt_5_590,.Wgt_5_591,.Wgt_5_592,.Wgt_5_593,.Wgt_5_594,.Wgt_5_595,.Wgt_5_596,.Wgt_5_597,.Wgt_5_598,.Wgt_5_599,.Wgt_5_600,.Wgt_5_601,.Wgt_5_602,.Wgt_5_603,.Wgt_5_604,.Wgt_5_605,.Wgt_5_606,.Wgt_5_607,.Wgt_5_608,.Wgt_5_609,.Wgt_5_610,.Wgt_5_611,.Wgt_5_612,.Wgt_5_613,.Wgt_5_614,.Wgt_5_615,.Wgt_5_616,.Wgt_5_617,.Wgt_5_618,.Wgt_5_619,.Wgt_5_620,.Wgt_5_621,.Wgt_5_622,.Wgt_5_623,.Wgt_5_624,.Wgt_5_625,.Wgt_5_626,.Wgt_5_627,.Wgt_5_628,.Wgt_5_629,.Wgt_5_630,.Wgt_5_631,.Wgt_5_632,.Wgt_5_633,.Wgt_5_634,.Wgt_5_635,.Wgt_5_636,.Wgt_5_637,.Wgt_5_638,.Wgt_5_639,.Wgt_5_640,.Wgt_5_641,.Wgt_5_642,.Wgt_5_643,.Wgt_5_644,.Wgt_5_645,.Wgt_5_646,.Wgt_5_647,.Wgt_5_648,.Wgt_5_649,.Wgt_5_650,.Wgt_5_651,.Wgt_5_652,.Wgt_5_653,.Wgt_5_654,.Wgt_5_655,.Wgt_5_656,.Wgt_5_657,.Wgt_5_658,.Wgt_5_659,.Wgt_5_660,.Wgt_5_661,.Wgt_5_662,.Wgt_5_663,.Wgt_5_664,.Wgt_5_665,.Wgt_5_666,.Wgt_5_667,.Wgt_5_668,.Wgt_5_669,.Wgt_5_670,.Wgt_5_671,.Wgt_5_672,.Wgt_5_673,.Wgt_5_674,.Wgt_5_675,.Wgt_5_676,.Wgt_5_677,.Wgt_5_678,.Wgt_5_679,.Wgt_5_680,.Wgt_5_681,.Wgt_5_682,.Wgt_5_683,.Wgt_5_684,.Wgt_5_685,.Wgt_5_686,.Wgt_5_687,.Wgt_5_688,.Wgt_5_689,.Wgt_5_690,.Wgt_5_691,.Wgt_5_692,.Wgt_5_693,.Wgt_5_694,.Wgt_5_695,.Wgt_5_696,.Wgt_5_697,.Wgt_5_698,.Wgt_5_699,.Wgt_5_700,.Wgt_5_701,.Wgt_5_702,.Wgt_5_703,.Wgt_5_704,.Wgt_5_705,.Wgt_5_706,.Wgt_5_707,.Wgt_5_708,.Wgt_5_709,.Wgt_5_710,.Wgt_5_711,.Wgt_5_712,.Wgt_5_713,.Wgt_5_714,.Wgt_5_715,.Wgt_5_716,.Wgt_5_717,.Wgt_5_718,.Wgt_5_719,.Wgt_5_720,.Wgt_5_721,.Wgt_5_722,.Wgt_5_723,.Wgt_5_724,.Wgt_5_725,.Wgt_5_726,.Wgt_5_727,.Wgt_5_728,.Wgt_5_729,.Wgt_5_730,.Wgt_5_731,.Wgt_5_732,.Wgt_5_733,.Wgt_5_734,.Wgt_5_735,.Wgt_5_736,.Wgt_5_737,.Wgt_5_738,.Wgt_5_739,.Wgt_5_740,.Wgt_5_741,.Wgt_5_742,.Wgt_5_743,.Wgt_5_744,.Wgt_5_745,.Wgt_5_746,.Wgt_5_747,.Wgt_5_748,.Wgt_5_749,.Wgt_5_750,.Wgt_5_751,.Wgt_5_752,.Wgt_5_753,.Wgt_5_754,.Wgt_5_755,.Wgt_5_756,.Wgt_5_757,.Wgt_5_758,.Wgt_5_759,.Wgt_5_760,.Wgt_5_761,.Wgt_5_762,.Wgt_5_763,.Wgt_5_764,.Wgt_5_765,.Wgt_5_766,.Wgt_5_767,.Wgt_5_768,.Wgt_5_769,.Wgt_5_770,.Wgt_5_771,.Wgt_5_772,.Wgt_5_773,.Wgt_5_774,.Wgt_5_775,.Wgt_5_776,.Wgt_5_777,.Wgt_5_778,.Wgt_5_779,.Wgt_5_780,.Wgt_5_781,.Wgt_5_782,.Wgt_5_783,.Wgt_5_784,
.Wgt_6_0,.Wgt_6_1,.Wgt_6_2,.Wgt_6_3,.Wgt_6_4,.Wgt_6_5,.Wgt_6_6,.Wgt_6_7,.Wgt_6_8,.Wgt_6_9,.Wgt_6_10,.Wgt_6_11,.Wgt_6_12,.Wgt_6_13,.Wgt_6_14,.Wgt_6_15,.Wgt_6_16,.Wgt_6_17,.Wgt_6_18,.Wgt_6_19,.Wgt_6_20,.Wgt_6_21,.Wgt_6_22,.Wgt_6_23,.Wgt_6_24,.Wgt_6_25,.Wgt_6_26,.Wgt_6_27,.Wgt_6_28,.Wgt_6_29,.Wgt_6_30,.Wgt_6_31,.Wgt_6_32,.Wgt_6_33,.Wgt_6_34,.Wgt_6_35,.Wgt_6_36,.Wgt_6_37,.Wgt_6_38,.Wgt_6_39,.Wgt_6_40,.Wgt_6_41,.Wgt_6_42,.Wgt_6_43,.Wgt_6_44,.Wgt_6_45,.Wgt_6_46,.Wgt_6_47,.Wgt_6_48,.Wgt_6_49,.Wgt_6_50,.Wgt_6_51,.Wgt_6_52,.Wgt_6_53,.Wgt_6_54,.Wgt_6_55,.Wgt_6_56,.Wgt_6_57,.Wgt_6_58,.Wgt_6_59,.Wgt_6_60,.Wgt_6_61,.Wgt_6_62,.Wgt_6_63,.Wgt_6_64,.Wgt_6_65,.Wgt_6_66,.Wgt_6_67,.Wgt_6_68,.Wgt_6_69,.Wgt_6_70,.Wgt_6_71,.Wgt_6_72,.Wgt_6_73,.Wgt_6_74,.Wgt_6_75,.Wgt_6_76,.Wgt_6_77,.Wgt_6_78,.Wgt_6_79,.Wgt_6_80,.Wgt_6_81,.Wgt_6_82,.Wgt_6_83,.Wgt_6_84,.Wgt_6_85,.Wgt_6_86,.Wgt_6_87,.Wgt_6_88,.Wgt_6_89,.Wgt_6_90,.Wgt_6_91,.Wgt_6_92,.Wgt_6_93,.Wgt_6_94,.Wgt_6_95,.Wgt_6_96,.Wgt_6_97,.Wgt_6_98,.Wgt_6_99,.Wgt_6_100,.Wgt_6_101,.Wgt_6_102,.Wgt_6_103,.Wgt_6_104,.Wgt_6_105,.Wgt_6_106,.Wgt_6_107,.Wgt_6_108,.Wgt_6_109,.Wgt_6_110,.Wgt_6_111,.Wgt_6_112,.Wgt_6_113,.Wgt_6_114,.Wgt_6_115,.Wgt_6_116,.Wgt_6_117,.Wgt_6_118,.Wgt_6_119,.Wgt_6_120,.Wgt_6_121,.Wgt_6_122,.Wgt_6_123,.Wgt_6_124,.Wgt_6_125,.Wgt_6_126,.Wgt_6_127,.Wgt_6_128,.Wgt_6_129,.Wgt_6_130,.Wgt_6_131,.Wgt_6_132,.Wgt_6_133,.Wgt_6_134,.Wgt_6_135,.Wgt_6_136,.Wgt_6_137,.Wgt_6_138,.Wgt_6_139,.Wgt_6_140,.Wgt_6_141,.Wgt_6_142,.Wgt_6_143,.Wgt_6_144,.Wgt_6_145,.Wgt_6_146,.Wgt_6_147,.Wgt_6_148,.Wgt_6_149,.Wgt_6_150,.Wgt_6_151,.Wgt_6_152,.Wgt_6_153,.Wgt_6_154,.Wgt_6_155,.Wgt_6_156,.Wgt_6_157,.Wgt_6_158,.Wgt_6_159,.Wgt_6_160,.Wgt_6_161,.Wgt_6_162,.Wgt_6_163,.Wgt_6_164,.Wgt_6_165,.Wgt_6_166,.Wgt_6_167,.Wgt_6_168,.Wgt_6_169,.Wgt_6_170,.Wgt_6_171,.Wgt_6_172,.Wgt_6_173,.Wgt_6_174,.Wgt_6_175,.Wgt_6_176,.Wgt_6_177,.Wgt_6_178,.Wgt_6_179,.Wgt_6_180,.Wgt_6_181,.Wgt_6_182,.Wgt_6_183,.Wgt_6_184,.Wgt_6_185,.Wgt_6_186,.Wgt_6_187,.Wgt_6_188,.Wgt_6_189,.Wgt_6_190,.Wgt_6_191,.Wgt_6_192,.Wgt_6_193,.Wgt_6_194,.Wgt_6_195,.Wgt_6_196,.Wgt_6_197,.Wgt_6_198,.Wgt_6_199,.Wgt_6_200,.Wgt_6_201,.Wgt_6_202,.Wgt_6_203,.Wgt_6_204,.Wgt_6_205,.Wgt_6_206,.Wgt_6_207,.Wgt_6_208,.Wgt_6_209,.Wgt_6_210,.Wgt_6_211,.Wgt_6_212,.Wgt_6_213,.Wgt_6_214,.Wgt_6_215,.Wgt_6_216,.Wgt_6_217,.Wgt_6_218,.Wgt_6_219,.Wgt_6_220,.Wgt_6_221,.Wgt_6_222,.Wgt_6_223,.Wgt_6_224,.Wgt_6_225,.Wgt_6_226,.Wgt_6_227,.Wgt_6_228,.Wgt_6_229,.Wgt_6_230,.Wgt_6_231,.Wgt_6_232,.Wgt_6_233,.Wgt_6_234,.Wgt_6_235,.Wgt_6_236,.Wgt_6_237,.Wgt_6_238,.Wgt_6_239,.Wgt_6_240,.Wgt_6_241,.Wgt_6_242,.Wgt_6_243,.Wgt_6_244,.Wgt_6_245,.Wgt_6_246,.Wgt_6_247,.Wgt_6_248,.Wgt_6_249,.Wgt_6_250,.Wgt_6_251,.Wgt_6_252,.Wgt_6_253,.Wgt_6_254,.Wgt_6_255,.Wgt_6_256,.Wgt_6_257,.Wgt_6_258,.Wgt_6_259,.Wgt_6_260,.Wgt_6_261,.Wgt_6_262,.Wgt_6_263,.Wgt_6_264,.Wgt_6_265,.Wgt_6_266,.Wgt_6_267,.Wgt_6_268,.Wgt_6_269,.Wgt_6_270,.Wgt_6_271,.Wgt_6_272,.Wgt_6_273,.Wgt_6_274,.Wgt_6_275,.Wgt_6_276,.Wgt_6_277,.Wgt_6_278,.Wgt_6_279,.Wgt_6_280,.Wgt_6_281,.Wgt_6_282,.Wgt_6_283,.Wgt_6_284,.Wgt_6_285,.Wgt_6_286,.Wgt_6_287,.Wgt_6_288,.Wgt_6_289,.Wgt_6_290,.Wgt_6_291,.Wgt_6_292,.Wgt_6_293,.Wgt_6_294,.Wgt_6_295,.Wgt_6_296,.Wgt_6_297,.Wgt_6_298,.Wgt_6_299,.Wgt_6_300,.Wgt_6_301,.Wgt_6_302,.Wgt_6_303,.Wgt_6_304,.Wgt_6_305,.Wgt_6_306,.Wgt_6_307,.Wgt_6_308,.Wgt_6_309,.Wgt_6_310,.Wgt_6_311,.Wgt_6_312,.Wgt_6_313,.Wgt_6_314,.Wgt_6_315,.Wgt_6_316,.Wgt_6_317,.Wgt_6_318,.Wgt_6_319,.Wgt_6_320,.Wgt_6_321,.Wgt_6_322,.Wgt_6_323,.Wgt_6_324,.Wgt_6_325,.Wgt_6_326,.Wgt_6_327,.Wgt_6_328,.Wgt_6_329,.Wgt_6_330,.Wgt_6_331,.Wgt_6_332,.Wgt_6_333,.Wgt_6_334,.Wgt_6_335,.Wgt_6_336,.Wgt_6_337,.Wgt_6_338,.Wgt_6_339,.Wgt_6_340,.Wgt_6_341,.Wgt_6_342,.Wgt_6_343,.Wgt_6_344,.Wgt_6_345,.Wgt_6_346,.Wgt_6_347,.Wgt_6_348,.Wgt_6_349,.Wgt_6_350,.Wgt_6_351,.Wgt_6_352,.Wgt_6_353,.Wgt_6_354,.Wgt_6_355,.Wgt_6_356,.Wgt_6_357,.Wgt_6_358,.Wgt_6_359,.Wgt_6_360,.Wgt_6_361,.Wgt_6_362,.Wgt_6_363,.Wgt_6_364,.Wgt_6_365,.Wgt_6_366,.Wgt_6_367,.Wgt_6_368,.Wgt_6_369,.Wgt_6_370,.Wgt_6_371,.Wgt_6_372,.Wgt_6_373,.Wgt_6_374,.Wgt_6_375,.Wgt_6_376,.Wgt_6_377,.Wgt_6_378,.Wgt_6_379,.Wgt_6_380,.Wgt_6_381,.Wgt_6_382,.Wgt_6_383,.Wgt_6_384,.Wgt_6_385,.Wgt_6_386,.Wgt_6_387,.Wgt_6_388,.Wgt_6_389,.Wgt_6_390,.Wgt_6_391,.Wgt_6_392,.Wgt_6_393,.Wgt_6_394,.Wgt_6_395,.Wgt_6_396,.Wgt_6_397,.Wgt_6_398,.Wgt_6_399,.Wgt_6_400,.Wgt_6_401,.Wgt_6_402,.Wgt_6_403,.Wgt_6_404,.Wgt_6_405,.Wgt_6_406,.Wgt_6_407,.Wgt_6_408,.Wgt_6_409,.Wgt_6_410,.Wgt_6_411,.Wgt_6_412,.Wgt_6_413,.Wgt_6_414,.Wgt_6_415,.Wgt_6_416,.Wgt_6_417,.Wgt_6_418,.Wgt_6_419,.Wgt_6_420,.Wgt_6_421,.Wgt_6_422,.Wgt_6_423,.Wgt_6_424,.Wgt_6_425,.Wgt_6_426,.Wgt_6_427,.Wgt_6_428,.Wgt_6_429,.Wgt_6_430,.Wgt_6_431,.Wgt_6_432,.Wgt_6_433,.Wgt_6_434,.Wgt_6_435,.Wgt_6_436,.Wgt_6_437,.Wgt_6_438,.Wgt_6_439,.Wgt_6_440,.Wgt_6_441,.Wgt_6_442,.Wgt_6_443,.Wgt_6_444,.Wgt_6_445,.Wgt_6_446,.Wgt_6_447,.Wgt_6_448,.Wgt_6_449,.Wgt_6_450,.Wgt_6_451,.Wgt_6_452,.Wgt_6_453,.Wgt_6_454,.Wgt_6_455,.Wgt_6_456,.Wgt_6_457,.Wgt_6_458,.Wgt_6_459,.Wgt_6_460,.Wgt_6_461,.Wgt_6_462,.Wgt_6_463,.Wgt_6_464,.Wgt_6_465,.Wgt_6_466,.Wgt_6_467,.Wgt_6_468,.Wgt_6_469,.Wgt_6_470,.Wgt_6_471,.Wgt_6_472,.Wgt_6_473,.Wgt_6_474,.Wgt_6_475,.Wgt_6_476,.Wgt_6_477,.Wgt_6_478,.Wgt_6_479,.Wgt_6_480,.Wgt_6_481,.Wgt_6_482,.Wgt_6_483,.Wgt_6_484,.Wgt_6_485,.Wgt_6_486,.Wgt_6_487,.Wgt_6_488,.Wgt_6_489,.Wgt_6_490,.Wgt_6_491,.Wgt_6_492,.Wgt_6_493,.Wgt_6_494,.Wgt_6_495,.Wgt_6_496,.Wgt_6_497,.Wgt_6_498,.Wgt_6_499,.Wgt_6_500,.Wgt_6_501,.Wgt_6_502,.Wgt_6_503,.Wgt_6_504,.Wgt_6_505,.Wgt_6_506,.Wgt_6_507,.Wgt_6_508,.Wgt_6_509,.Wgt_6_510,.Wgt_6_511,.Wgt_6_512,.Wgt_6_513,.Wgt_6_514,.Wgt_6_515,.Wgt_6_516,.Wgt_6_517,.Wgt_6_518,.Wgt_6_519,.Wgt_6_520,.Wgt_6_521,.Wgt_6_522,.Wgt_6_523,.Wgt_6_524,.Wgt_6_525,.Wgt_6_526,.Wgt_6_527,.Wgt_6_528,.Wgt_6_529,.Wgt_6_530,.Wgt_6_531,.Wgt_6_532,.Wgt_6_533,.Wgt_6_534,.Wgt_6_535,.Wgt_6_536,.Wgt_6_537,.Wgt_6_538,.Wgt_6_539,.Wgt_6_540,.Wgt_6_541,.Wgt_6_542,.Wgt_6_543,.Wgt_6_544,.Wgt_6_545,.Wgt_6_546,.Wgt_6_547,.Wgt_6_548,.Wgt_6_549,.Wgt_6_550,.Wgt_6_551,.Wgt_6_552,.Wgt_6_553,.Wgt_6_554,.Wgt_6_555,.Wgt_6_556,.Wgt_6_557,.Wgt_6_558,.Wgt_6_559,.Wgt_6_560,.Wgt_6_561,.Wgt_6_562,.Wgt_6_563,.Wgt_6_564,.Wgt_6_565,.Wgt_6_566,.Wgt_6_567,.Wgt_6_568,.Wgt_6_569,.Wgt_6_570,.Wgt_6_571,.Wgt_6_572,.Wgt_6_573,.Wgt_6_574,.Wgt_6_575,.Wgt_6_576,.Wgt_6_577,.Wgt_6_578,.Wgt_6_579,.Wgt_6_580,.Wgt_6_581,.Wgt_6_582,.Wgt_6_583,.Wgt_6_584,.Wgt_6_585,.Wgt_6_586,.Wgt_6_587,.Wgt_6_588,.Wgt_6_589,.Wgt_6_590,.Wgt_6_591,.Wgt_6_592,.Wgt_6_593,.Wgt_6_594,.Wgt_6_595,.Wgt_6_596,.Wgt_6_597,.Wgt_6_598,.Wgt_6_599,.Wgt_6_600,.Wgt_6_601,.Wgt_6_602,.Wgt_6_603,.Wgt_6_604,.Wgt_6_605,.Wgt_6_606,.Wgt_6_607,.Wgt_6_608,.Wgt_6_609,.Wgt_6_610,.Wgt_6_611,.Wgt_6_612,.Wgt_6_613,.Wgt_6_614,.Wgt_6_615,.Wgt_6_616,.Wgt_6_617,.Wgt_6_618,.Wgt_6_619,.Wgt_6_620,.Wgt_6_621,.Wgt_6_622,.Wgt_6_623,.Wgt_6_624,.Wgt_6_625,.Wgt_6_626,.Wgt_6_627,.Wgt_6_628,.Wgt_6_629,.Wgt_6_630,.Wgt_6_631,.Wgt_6_632,.Wgt_6_633,.Wgt_6_634,.Wgt_6_635,.Wgt_6_636,.Wgt_6_637,.Wgt_6_638,.Wgt_6_639,.Wgt_6_640,.Wgt_6_641,.Wgt_6_642,.Wgt_6_643,.Wgt_6_644,.Wgt_6_645,.Wgt_6_646,.Wgt_6_647,.Wgt_6_648,.Wgt_6_649,.Wgt_6_650,.Wgt_6_651,.Wgt_6_652,.Wgt_6_653,.Wgt_6_654,.Wgt_6_655,.Wgt_6_656,.Wgt_6_657,.Wgt_6_658,.Wgt_6_659,.Wgt_6_660,.Wgt_6_661,.Wgt_6_662,.Wgt_6_663,.Wgt_6_664,.Wgt_6_665,.Wgt_6_666,.Wgt_6_667,.Wgt_6_668,.Wgt_6_669,.Wgt_6_670,.Wgt_6_671,.Wgt_6_672,.Wgt_6_673,.Wgt_6_674,.Wgt_6_675,.Wgt_6_676,.Wgt_6_677,.Wgt_6_678,.Wgt_6_679,.Wgt_6_680,.Wgt_6_681,.Wgt_6_682,.Wgt_6_683,.Wgt_6_684,.Wgt_6_685,.Wgt_6_686,.Wgt_6_687,.Wgt_6_688,.Wgt_6_689,.Wgt_6_690,.Wgt_6_691,.Wgt_6_692,.Wgt_6_693,.Wgt_6_694,.Wgt_6_695,.Wgt_6_696,.Wgt_6_697,.Wgt_6_698,.Wgt_6_699,.Wgt_6_700,.Wgt_6_701,.Wgt_6_702,.Wgt_6_703,.Wgt_6_704,.Wgt_6_705,.Wgt_6_706,.Wgt_6_707,.Wgt_6_708,.Wgt_6_709,.Wgt_6_710,.Wgt_6_711,.Wgt_6_712,.Wgt_6_713,.Wgt_6_714,.Wgt_6_715,.Wgt_6_716,.Wgt_6_717,.Wgt_6_718,.Wgt_6_719,.Wgt_6_720,.Wgt_6_721,.Wgt_6_722,.Wgt_6_723,.Wgt_6_724,.Wgt_6_725,.Wgt_6_726,.Wgt_6_727,.Wgt_6_728,.Wgt_6_729,.Wgt_6_730,.Wgt_6_731,.Wgt_6_732,.Wgt_6_733,.Wgt_6_734,.Wgt_6_735,.Wgt_6_736,.Wgt_6_737,.Wgt_6_738,.Wgt_6_739,.Wgt_6_740,.Wgt_6_741,.Wgt_6_742,.Wgt_6_743,.Wgt_6_744,.Wgt_6_745,.Wgt_6_746,.Wgt_6_747,.Wgt_6_748,.Wgt_6_749,.Wgt_6_750,.Wgt_6_751,.Wgt_6_752,.Wgt_6_753,.Wgt_6_754,.Wgt_6_755,.Wgt_6_756,.Wgt_6_757,.Wgt_6_758,.Wgt_6_759,.Wgt_6_760,.Wgt_6_761,.Wgt_6_762,.Wgt_6_763,.Wgt_6_764,.Wgt_6_765,.Wgt_6_766,.Wgt_6_767,.Wgt_6_768,.Wgt_6_769,.Wgt_6_770,.Wgt_6_771,.Wgt_6_772,.Wgt_6_773,.Wgt_6_774,.Wgt_6_775,.Wgt_6_776,.Wgt_6_777,.Wgt_6_778,.Wgt_6_779,.Wgt_6_780,.Wgt_6_781,.Wgt_6_782,.Wgt_6_783,.Wgt_6_784,
.Wgt_7_0,.Wgt_7_1,.Wgt_7_2,.Wgt_7_3,.Wgt_7_4,.Wgt_7_5,.Wgt_7_6,.Wgt_7_7,.Wgt_7_8,.Wgt_7_9,.Wgt_7_10,.Wgt_7_11,.Wgt_7_12,.Wgt_7_13,.Wgt_7_14,.Wgt_7_15,.Wgt_7_16,.Wgt_7_17,.Wgt_7_18,.Wgt_7_19,.Wgt_7_20,.Wgt_7_21,.Wgt_7_22,.Wgt_7_23,.Wgt_7_24,.Wgt_7_25,.Wgt_7_26,.Wgt_7_27,.Wgt_7_28,.Wgt_7_29,.Wgt_7_30,.Wgt_7_31,.Wgt_7_32,.Wgt_7_33,.Wgt_7_34,.Wgt_7_35,.Wgt_7_36,.Wgt_7_37,.Wgt_7_38,.Wgt_7_39,.Wgt_7_40,.Wgt_7_41,.Wgt_7_42,.Wgt_7_43,.Wgt_7_44,.Wgt_7_45,.Wgt_7_46,.Wgt_7_47,.Wgt_7_48,.Wgt_7_49,.Wgt_7_50,.Wgt_7_51,.Wgt_7_52,.Wgt_7_53,.Wgt_7_54,.Wgt_7_55,.Wgt_7_56,.Wgt_7_57,.Wgt_7_58,.Wgt_7_59,.Wgt_7_60,.Wgt_7_61,.Wgt_7_62,.Wgt_7_63,.Wgt_7_64,.Wgt_7_65,.Wgt_7_66,.Wgt_7_67,.Wgt_7_68,.Wgt_7_69,.Wgt_7_70,.Wgt_7_71,.Wgt_7_72,.Wgt_7_73,.Wgt_7_74,.Wgt_7_75,.Wgt_7_76,.Wgt_7_77,.Wgt_7_78,.Wgt_7_79,.Wgt_7_80,.Wgt_7_81,.Wgt_7_82,.Wgt_7_83,.Wgt_7_84,.Wgt_7_85,.Wgt_7_86,.Wgt_7_87,.Wgt_7_88,.Wgt_7_89,.Wgt_7_90,.Wgt_7_91,.Wgt_7_92,.Wgt_7_93,.Wgt_7_94,.Wgt_7_95,.Wgt_7_96,.Wgt_7_97,.Wgt_7_98,.Wgt_7_99,.Wgt_7_100,.Wgt_7_101,.Wgt_7_102,.Wgt_7_103,.Wgt_7_104,.Wgt_7_105,.Wgt_7_106,.Wgt_7_107,.Wgt_7_108,.Wgt_7_109,.Wgt_7_110,.Wgt_7_111,.Wgt_7_112,.Wgt_7_113,.Wgt_7_114,.Wgt_7_115,.Wgt_7_116,.Wgt_7_117,.Wgt_7_118,.Wgt_7_119,.Wgt_7_120,.Wgt_7_121,.Wgt_7_122,.Wgt_7_123,.Wgt_7_124,.Wgt_7_125,.Wgt_7_126,.Wgt_7_127,.Wgt_7_128,.Wgt_7_129,.Wgt_7_130,.Wgt_7_131,.Wgt_7_132,.Wgt_7_133,.Wgt_7_134,.Wgt_7_135,.Wgt_7_136,.Wgt_7_137,.Wgt_7_138,.Wgt_7_139,.Wgt_7_140,.Wgt_7_141,.Wgt_7_142,.Wgt_7_143,.Wgt_7_144,.Wgt_7_145,.Wgt_7_146,.Wgt_7_147,.Wgt_7_148,.Wgt_7_149,.Wgt_7_150,.Wgt_7_151,.Wgt_7_152,.Wgt_7_153,.Wgt_7_154,.Wgt_7_155,.Wgt_7_156,.Wgt_7_157,.Wgt_7_158,.Wgt_7_159,.Wgt_7_160,.Wgt_7_161,.Wgt_7_162,.Wgt_7_163,.Wgt_7_164,.Wgt_7_165,.Wgt_7_166,.Wgt_7_167,.Wgt_7_168,.Wgt_7_169,.Wgt_7_170,.Wgt_7_171,.Wgt_7_172,.Wgt_7_173,.Wgt_7_174,.Wgt_7_175,.Wgt_7_176,.Wgt_7_177,.Wgt_7_178,.Wgt_7_179,.Wgt_7_180,.Wgt_7_181,.Wgt_7_182,.Wgt_7_183,.Wgt_7_184,.Wgt_7_185,.Wgt_7_186,.Wgt_7_187,.Wgt_7_188,.Wgt_7_189,.Wgt_7_190,.Wgt_7_191,.Wgt_7_192,.Wgt_7_193,.Wgt_7_194,.Wgt_7_195,.Wgt_7_196,.Wgt_7_197,.Wgt_7_198,.Wgt_7_199,.Wgt_7_200,.Wgt_7_201,.Wgt_7_202,.Wgt_7_203,.Wgt_7_204,.Wgt_7_205,.Wgt_7_206,.Wgt_7_207,.Wgt_7_208,.Wgt_7_209,.Wgt_7_210,.Wgt_7_211,.Wgt_7_212,.Wgt_7_213,.Wgt_7_214,.Wgt_7_215,.Wgt_7_216,.Wgt_7_217,.Wgt_7_218,.Wgt_7_219,.Wgt_7_220,.Wgt_7_221,.Wgt_7_222,.Wgt_7_223,.Wgt_7_224,.Wgt_7_225,.Wgt_7_226,.Wgt_7_227,.Wgt_7_228,.Wgt_7_229,.Wgt_7_230,.Wgt_7_231,.Wgt_7_232,.Wgt_7_233,.Wgt_7_234,.Wgt_7_235,.Wgt_7_236,.Wgt_7_237,.Wgt_7_238,.Wgt_7_239,.Wgt_7_240,.Wgt_7_241,.Wgt_7_242,.Wgt_7_243,.Wgt_7_244,.Wgt_7_245,.Wgt_7_246,.Wgt_7_247,.Wgt_7_248,.Wgt_7_249,.Wgt_7_250,.Wgt_7_251,.Wgt_7_252,.Wgt_7_253,.Wgt_7_254,.Wgt_7_255,.Wgt_7_256,.Wgt_7_257,.Wgt_7_258,.Wgt_7_259,.Wgt_7_260,.Wgt_7_261,.Wgt_7_262,.Wgt_7_263,.Wgt_7_264,.Wgt_7_265,.Wgt_7_266,.Wgt_7_267,.Wgt_7_268,.Wgt_7_269,.Wgt_7_270,.Wgt_7_271,.Wgt_7_272,.Wgt_7_273,.Wgt_7_274,.Wgt_7_275,.Wgt_7_276,.Wgt_7_277,.Wgt_7_278,.Wgt_7_279,.Wgt_7_280,.Wgt_7_281,.Wgt_7_282,.Wgt_7_283,.Wgt_7_284,.Wgt_7_285,.Wgt_7_286,.Wgt_7_287,.Wgt_7_288,.Wgt_7_289,.Wgt_7_290,.Wgt_7_291,.Wgt_7_292,.Wgt_7_293,.Wgt_7_294,.Wgt_7_295,.Wgt_7_296,.Wgt_7_297,.Wgt_7_298,.Wgt_7_299,.Wgt_7_300,.Wgt_7_301,.Wgt_7_302,.Wgt_7_303,.Wgt_7_304,.Wgt_7_305,.Wgt_7_306,.Wgt_7_307,.Wgt_7_308,.Wgt_7_309,.Wgt_7_310,.Wgt_7_311,.Wgt_7_312,.Wgt_7_313,.Wgt_7_314,.Wgt_7_315,.Wgt_7_316,.Wgt_7_317,.Wgt_7_318,.Wgt_7_319,.Wgt_7_320,.Wgt_7_321,.Wgt_7_322,.Wgt_7_323,.Wgt_7_324,.Wgt_7_325,.Wgt_7_326,.Wgt_7_327,.Wgt_7_328,.Wgt_7_329,.Wgt_7_330,.Wgt_7_331,.Wgt_7_332,.Wgt_7_333,.Wgt_7_334,.Wgt_7_335,.Wgt_7_336,.Wgt_7_337,.Wgt_7_338,.Wgt_7_339,.Wgt_7_340,.Wgt_7_341,.Wgt_7_342,.Wgt_7_343,.Wgt_7_344,.Wgt_7_345,.Wgt_7_346,.Wgt_7_347,.Wgt_7_348,.Wgt_7_349,.Wgt_7_350,.Wgt_7_351,.Wgt_7_352,.Wgt_7_353,.Wgt_7_354,.Wgt_7_355,.Wgt_7_356,.Wgt_7_357,.Wgt_7_358,.Wgt_7_359,.Wgt_7_360,.Wgt_7_361,.Wgt_7_362,.Wgt_7_363,.Wgt_7_364,.Wgt_7_365,.Wgt_7_366,.Wgt_7_367,.Wgt_7_368,.Wgt_7_369,.Wgt_7_370,.Wgt_7_371,.Wgt_7_372,.Wgt_7_373,.Wgt_7_374,.Wgt_7_375,.Wgt_7_376,.Wgt_7_377,.Wgt_7_378,.Wgt_7_379,.Wgt_7_380,.Wgt_7_381,.Wgt_7_382,.Wgt_7_383,.Wgt_7_384,.Wgt_7_385,.Wgt_7_386,.Wgt_7_387,.Wgt_7_388,.Wgt_7_389,.Wgt_7_390,.Wgt_7_391,.Wgt_7_392,.Wgt_7_393,.Wgt_7_394,.Wgt_7_395,.Wgt_7_396,.Wgt_7_397,.Wgt_7_398,.Wgt_7_399,.Wgt_7_400,.Wgt_7_401,.Wgt_7_402,.Wgt_7_403,.Wgt_7_404,.Wgt_7_405,.Wgt_7_406,.Wgt_7_407,.Wgt_7_408,.Wgt_7_409,.Wgt_7_410,.Wgt_7_411,.Wgt_7_412,.Wgt_7_413,.Wgt_7_414,.Wgt_7_415,.Wgt_7_416,.Wgt_7_417,.Wgt_7_418,.Wgt_7_419,.Wgt_7_420,.Wgt_7_421,.Wgt_7_422,.Wgt_7_423,.Wgt_7_424,.Wgt_7_425,.Wgt_7_426,.Wgt_7_427,.Wgt_7_428,.Wgt_7_429,.Wgt_7_430,.Wgt_7_431,.Wgt_7_432,.Wgt_7_433,.Wgt_7_434,.Wgt_7_435,.Wgt_7_436,.Wgt_7_437,.Wgt_7_438,.Wgt_7_439,.Wgt_7_440,.Wgt_7_441,.Wgt_7_442,.Wgt_7_443,.Wgt_7_444,.Wgt_7_445,.Wgt_7_446,.Wgt_7_447,.Wgt_7_448,.Wgt_7_449,.Wgt_7_450,.Wgt_7_451,.Wgt_7_452,.Wgt_7_453,.Wgt_7_454,.Wgt_7_455,.Wgt_7_456,.Wgt_7_457,.Wgt_7_458,.Wgt_7_459,.Wgt_7_460,.Wgt_7_461,.Wgt_7_462,.Wgt_7_463,.Wgt_7_464,.Wgt_7_465,.Wgt_7_466,.Wgt_7_467,.Wgt_7_468,.Wgt_7_469,.Wgt_7_470,.Wgt_7_471,.Wgt_7_472,.Wgt_7_473,.Wgt_7_474,.Wgt_7_475,.Wgt_7_476,.Wgt_7_477,.Wgt_7_478,.Wgt_7_479,.Wgt_7_480,.Wgt_7_481,.Wgt_7_482,.Wgt_7_483,.Wgt_7_484,.Wgt_7_485,.Wgt_7_486,.Wgt_7_487,.Wgt_7_488,.Wgt_7_489,.Wgt_7_490,.Wgt_7_491,.Wgt_7_492,.Wgt_7_493,.Wgt_7_494,.Wgt_7_495,.Wgt_7_496,.Wgt_7_497,.Wgt_7_498,.Wgt_7_499,.Wgt_7_500,.Wgt_7_501,.Wgt_7_502,.Wgt_7_503,.Wgt_7_504,.Wgt_7_505,.Wgt_7_506,.Wgt_7_507,.Wgt_7_508,.Wgt_7_509,.Wgt_7_510,.Wgt_7_511,.Wgt_7_512,.Wgt_7_513,.Wgt_7_514,.Wgt_7_515,.Wgt_7_516,.Wgt_7_517,.Wgt_7_518,.Wgt_7_519,.Wgt_7_520,.Wgt_7_521,.Wgt_7_522,.Wgt_7_523,.Wgt_7_524,.Wgt_7_525,.Wgt_7_526,.Wgt_7_527,.Wgt_7_528,.Wgt_7_529,.Wgt_7_530,.Wgt_7_531,.Wgt_7_532,.Wgt_7_533,.Wgt_7_534,.Wgt_7_535,.Wgt_7_536,.Wgt_7_537,.Wgt_7_538,.Wgt_7_539,.Wgt_7_540,.Wgt_7_541,.Wgt_7_542,.Wgt_7_543,.Wgt_7_544,.Wgt_7_545,.Wgt_7_546,.Wgt_7_547,.Wgt_7_548,.Wgt_7_549,.Wgt_7_550,.Wgt_7_551,.Wgt_7_552,.Wgt_7_553,.Wgt_7_554,.Wgt_7_555,.Wgt_7_556,.Wgt_7_557,.Wgt_7_558,.Wgt_7_559,.Wgt_7_560,.Wgt_7_561,.Wgt_7_562,.Wgt_7_563,.Wgt_7_564,.Wgt_7_565,.Wgt_7_566,.Wgt_7_567,.Wgt_7_568,.Wgt_7_569,.Wgt_7_570,.Wgt_7_571,.Wgt_7_572,.Wgt_7_573,.Wgt_7_574,.Wgt_7_575,.Wgt_7_576,.Wgt_7_577,.Wgt_7_578,.Wgt_7_579,.Wgt_7_580,.Wgt_7_581,.Wgt_7_582,.Wgt_7_583,.Wgt_7_584,.Wgt_7_585,.Wgt_7_586,.Wgt_7_587,.Wgt_7_588,.Wgt_7_589,.Wgt_7_590,.Wgt_7_591,.Wgt_7_592,.Wgt_7_593,.Wgt_7_594,.Wgt_7_595,.Wgt_7_596,.Wgt_7_597,.Wgt_7_598,.Wgt_7_599,.Wgt_7_600,.Wgt_7_601,.Wgt_7_602,.Wgt_7_603,.Wgt_7_604,.Wgt_7_605,.Wgt_7_606,.Wgt_7_607,.Wgt_7_608,.Wgt_7_609,.Wgt_7_610,.Wgt_7_611,.Wgt_7_612,.Wgt_7_613,.Wgt_7_614,.Wgt_7_615,.Wgt_7_616,.Wgt_7_617,.Wgt_7_618,.Wgt_7_619,.Wgt_7_620,.Wgt_7_621,.Wgt_7_622,.Wgt_7_623,.Wgt_7_624,.Wgt_7_625,.Wgt_7_626,.Wgt_7_627,.Wgt_7_628,.Wgt_7_629,.Wgt_7_630,.Wgt_7_631,.Wgt_7_632,.Wgt_7_633,.Wgt_7_634,.Wgt_7_635,.Wgt_7_636,.Wgt_7_637,.Wgt_7_638,.Wgt_7_639,.Wgt_7_640,.Wgt_7_641,.Wgt_7_642,.Wgt_7_643,.Wgt_7_644,.Wgt_7_645,.Wgt_7_646,.Wgt_7_647,.Wgt_7_648,.Wgt_7_649,.Wgt_7_650,.Wgt_7_651,.Wgt_7_652,.Wgt_7_653,.Wgt_7_654,.Wgt_7_655,.Wgt_7_656,.Wgt_7_657,.Wgt_7_658,.Wgt_7_659,.Wgt_7_660,.Wgt_7_661,.Wgt_7_662,.Wgt_7_663,.Wgt_7_664,.Wgt_7_665,.Wgt_7_666,.Wgt_7_667,.Wgt_7_668,.Wgt_7_669,.Wgt_7_670,.Wgt_7_671,.Wgt_7_672,.Wgt_7_673,.Wgt_7_674,.Wgt_7_675,.Wgt_7_676,.Wgt_7_677,.Wgt_7_678,.Wgt_7_679,.Wgt_7_680,.Wgt_7_681,.Wgt_7_682,.Wgt_7_683,.Wgt_7_684,.Wgt_7_685,.Wgt_7_686,.Wgt_7_687,.Wgt_7_688,.Wgt_7_689,.Wgt_7_690,.Wgt_7_691,.Wgt_7_692,.Wgt_7_693,.Wgt_7_694,.Wgt_7_695,.Wgt_7_696,.Wgt_7_697,.Wgt_7_698,.Wgt_7_699,.Wgt_7_700,.Wgt_7_701,.Wgt_7_702,.Wgt_7_703,.Wgt_7_704,.Wgt_7_705,.Wgt_7_706,.Wgt_7_707,.Wgt_7_708,.Wgt_7_709,.Wgt_7_710,.Wgt_7_711,.Wgt_7_712,.Wgt_7_713,.Wgt_7_714,.Wgt_7_715,.Wgt_7_716,.Wgt_7_717,.Wgt_7_718,.Wgt_7_719,.Wgt_7_720,.Wgt_7_721,.Wgt_7_722,.Wgt_7_723,.Wgt_7_724,.Wgt_7_725,.Wgt_7_726,.Wgt_7_727,.Wgt_7_728,.Wgt_7_729,.Wgt_7_730,.Wgt_7_731,.Wgt_7_732,.Wgt_7_733,.Wgt_7_734,.Wgt_7_735,.Wgt_7_736,.Wgt_7_737,.Wgt_7_738,.Wgt_7_739,.Wgt_7_740,.Wgt_7_741,.Wgt_7_742,.Wgt_7_743,.Wgt_7_744,.Wgt_7_745,.Wgt_7_746,.Wgt_7_747,.Wgt_7_748,.Wgt_7_749,.Wgt_7_750,.Wgt_7_751,.Wgt_7_752,.Wgt_7_753,.Wgt_7_754,.Wgt_7_755,.Wgt_7_756,.Wgt_7_757,.Wgt_7_758,.Wgt_7_759,.Wgt_7_760,.Wgt_7_761,.Wgt_7_762,.Wgt_7_763,.Wgt_7_764,.Wgt_7_765,.Wgt_7_766,.Wgt_7_767,.Wgt_7_768,.Wgt_7_769,.Wgt_7_770,.Wgt_7_771,.Wgt_7_772,.Wgt_7_773,.Wgt_7_774,.Wgt_7_775,.Wgt_7_776,.Wgt_7_777,.Wgt_7_778,.Wgt_7_779,.Wgt_7_780,.Wgt_7_781,.Wgt_7_782,.Wgt_7_783,.Wgt_7_784,
.Wgt_8_0,.Wgt_8_1,.Wgt_8_2,.Wgt_8_3,.Wgt_8_4,.Wgt_8_5,.Wgt_8_6,.Wgt_8_7,.Wgt_8_8,.Wgt_8_9,.Wgt_8_10,.Wgt_8_11,.Wgt_8_12,.Wgt_8_13,.Wgt_8_14,.Wgt_8_15,.Wgt_8_16,.Wgt_8_17,.Wgt_8_18,.Wgt_8_19,.Wgt_8_20,.Wgt_8_21,.Wgt_8_22,.Wgt_8_23,.Wgt_8_24,.Wgt_8_25,.Wgt_8_26,.Wgt_8_27,.Wgt_8_28,.Wgt_8_29,.Wgt_8_30,.Wgt_8_31,.Wgt_8_32,.Wgt_8_33,.Wgt_8_34,.Wgt_8_35,.Wgt_8_36,.Wgt_8_37,.Wgt_8_38,.Wgt_8_39,.Wgt_8_40,.Wgt_8_41,.Wgt_8_42,.Wgt_8_43,.Wgt_8_44,.Wgt_8_45,.Wgt_8_46,.Wgt_8_47,.Wgt_8_48,.Wgt_8_49,.Wgt_8_50,.Wgt_8_51,.Wgt_8_52,.Wgt_8_53,.Wgt_8_54,.Wgt_8_55,.Wgt_8_56,.Wgt_8_57,.Wgt_8_58,.Wgt_8_59,.Wgt_8_60,.Wgt_8_61,.Wgt_8_62,.Wgt_8_63,.Wgt_8_64,.Wgt_8_65,.Wgt_8_66,.Wgt_8_67,.Wgt_8_68,.Wgt_8_69,.Wgt_8_70,.Wgt_8_71,.Wgt_8_72,.Wgt_8_73,.Wgt_8_74,.Wgt_8_75,.Wgt_8_76,.Wgt_8_77,.Wgt_8_78,.Wgt_8_79,.Wgt_8_80,.Wgt_8_81,.Wgt_8_82,.Wgt_8_83,.Wgt_8_84,.Wgt_8_85,.Wgt_8_86,.Wgt_8_87,.Wgt_8_88,.Wgt_8_89,.Wgt_8_90,.Wgt_8_91,.Wgt_8_92,.Wgt_8_93,.Wgt_8_94,.Wgt_8_95,.Wgt_8_96,.Wgt_8_97,.Wgt_8_98,.Wgt_8_99,.Wgt_8_100,.Wgt_8_101,.Wgt_8_102,.Wgt_8_103,.Wgt_8_104,.Wgt_8_105,.Wgt_8_106,.Wgt_8_107,.Wgt_8_108,.Wgt_8_109,.Wgt_8_110,.Wgt_8_111,.Wgt_8_112,.Wgt_8_113,.Wgt_8_114,.Wgt_8_115,.Wgt_8_116,.Wgt_8_117,.Wgt_8_118,.Wgt_8_119,.Wgt_8_120,.Wgt_8_121,.Wgt_8_122,.Wgt_8_123,.Wgt_8_124,.Wgt_8_125,.Wgt_8_126,.Wgt_8_127,.Wgt_8_128,.Wgt_8_129,.Wgt_8_130,.Wgt_8_131,.Wgt_8_132,.Wgt_8_133,.Wgt_8_134,.Wgt_8_135,.Wgt_8_136,.Wgt_8_137,.Wgt_8_138,.Wgt_8_139,.Wgt_8_140,.Wgt_8_141,.Wgt_8_142,.Wgt_8_143,.Wgt_8_144,.Wgt_8_145,.Wgt_8_146,.Wgt_8_147,.Wgt_8_148,.Wgt_8_149,.Wgt_8_150,.Wgt_8_151,.Wgt_8_152,.Wgt_8_153,.Wgt_8_154,.Wgt_8_155,.Wgt_8_156,.Wgt_8_157,.Wgt_8_158,.Wgt_8_159,.Wgt_8_160,.Wgt_8_161,.Wgt_8_162,.Wgt_8_163,.Wgt_8_164,.Wgt_8_165,.Wgt_8_166,.Wgt_8_167,.Wgt_8_168,.Wgt_8_169,.Wgt_8_170,.Wgt_8_171,.Wgt_8_172,.Wgt_8_173,.Wgt_8_174,.Wgt_8_175,.Wgt_8_176,.Wgt_8_177,.Wgt_8_178,.Wgt_8_179,.Wgt_8_180,.Wgt_8_181,.Wgt_8_182,.Wgt_8_183,.Wgt_8_184,.Wgt_8_185,.Wgt_8_186,.Wgt_8_187,.Wgt_8_188,.Wgt_8_189,.Wgt_8_190,.Wgt_8_191,.Wgt_8_192,.Wgt_8_193,.Wgt_8_194,.Wgt_8_195,.Wgt_8_196,.Wgt_8_197,.Wgt_8_198,.Wgt_8_199,.Wgt_8_200,.Wgt_8_201,.Wgt_8_202,.Wgt_8_203,.Wgt_8_204,.Wgt_8_205,.Wgt_8_206,.Wgt_8_207,.Wgt_8_208,.Wgt_8_209,.Wgt_8_210,.Wgt_8_211,.Wgt_8_212,.Wgt_8_213,.Wgt_8_214,.Wgt_8_215,.Wgt_8_216,.Wgt_8_217,.Wgt_8_218,.Wgt_8_219,.Wgt_8_220,.Wgt_8_221,.Wgt_8_222,.Wgt_8_223,.Wgt_8_224,.Wgt_8_225,.Wgt_8_226,.Wgt_8_227,.Wgt_8_228,.Wgt_8_229,.Wgt_8_230,.Wgt_8_231,.Wgt_8_232,.Wgt_8_233,.Wgt_8_234,.Wgt_8_235,.Wgt_8_236,.Wgt_8_237,.Wgt_8_238,.Wgt_8_239,.Wgt_8_240,.Wgt_8_241,.Wgt_8_242,.Wgt_8_243,.Wgt_8_244,.Wgt_8_245,.Wgt_8_246,.Wgt_8_247,.Wgt_8_248,.Wgt_8_249,.Wgt_8_250,.Wgt_8_251,.Wgt_8_252,.Wgt_8_253,.Wgt_8_254,.Wgt_8_255,.Wgt_8_256,.Wgt_8_257,.Wgt_8_258,.Wgt_8_259,.Wgt_8_260,.Wgt_8_261,.Wgt_8_262,.Wgt_8_263,.Wgt_8_264,.Wgt_8_265,.Wgt_8_266,.Wgt_8_267,.Wgt_8_268,.Wgt_8_269,.Wgt_8_270,.Wgt_8_271,.Wgt_8_272,.Wgt_8_273,.Wgt_8_274,.Wgt_8_275,.Wgt_8_276,.Wgt_8_277,.Wgt_8_278,.Wgt_8_279,.Wgt_8_280,.Wgt_8_281,.Wgt_8_282,.Wgt_8_283,.Wgt_8_284,.Wgt_8_285,.Wgt_8_286,.Wgt_8_287,.Wgt_8_288,.Wgt_8_289,.Wgt_8_290,.Wgt_8_291,.Wgt_8_292,.Wgt_8_293,.Wgt_8_294,.Wgt_8_295,.Wgt_8_296,.Wgt_8_297,.Wgt_8_298,.Wgt_8_299,.Wgt_8_300,.Wgt_8_301,.Wgt_8_302,.Wgt_8_303,.Wgt_8_304,.Wgt_8_305,.Wgt_8_306,.Wgt_8_307,.Wgt_8_308,.Wgt_8_309,.Wgt_8_310,.Wgt_8_311,.Wgt_8_312,.Wgt_8_313,.Wgt_8_314,.Wgt_8_315,.Wgt_8_316,.Wgt_8_317,.Wgt_8_318,.Wgt_8_319,.Wgt_8_320,.Wgt_8_321,.Wgt_8_322,.Wgt_8_323,.Wgt_8_324,.Wgt_8_325,.Wgt_8_326,.Wgt_8_327,.Wgt_8_328,.Wgt_8_329,.Wgt_8_330,.Wgt_8_331,.Wgt_8_332,.Wgt_8_333,.Wgt_8_334,.Wgt_8_335,.Wgt_8_336,.Wgt_8_337,.Wgt_8_338,.Wgt_8_339,.Wgt_8_340,.Wgt_8_341,.Wgt_8_342,.Wgt_8_343,.Wgt_8_344,.Wgt_8_345,.Wgt_8_346,.Wgt_8_347,.Wgt_8_348,.Wgt_8_349,.Wgt_8_350,.Wgt_8_351,.Wgt_8_352,.Wgt_8_353,.Wgt_8_354,.Wgt_8_355,.Wgt_8_356,.Wgt_8_357,.Wgt_8_358,.Wgt_8_359,.Wgt_8_360,.Wgt_8_361,.Wgt_8_362,.Wgt_8_363,.Wgt_8_364,.Wgt_8_365,.Wgt_8_366,.Wgt_8_367,.Wgt_8_368,.Wgt_8_369,.Wgt_8_370,.Wgt_8_371,.Wgt_8_372,.Wgt_8_373,.Wgt_8_374,.Wgt_8_375,.Wgt_8_376,.Wgt_8_377,.Wgt_8_378,.Wgt_8_379,.Wgt_8_380,.Wgt_8_381,.Wgt_8_382,.Wgt_8_383,.Wgt_8_384,.Wgt_8_385,.Wgt_8_386,.Wgt_8_387,.Wgt_8_388,.Wgt_8_389,.Wgt_8_390,.Wgt_8_391,.Wgt_8_392,.Wgt_8_393,.Wgt_8_394,.Wgt_8_395,.Wgt_8_396,.Wgt_8_397,.Wgt_8_398,.Wgt_8_399,.Wgt_8_400,.Wgt_8_401,.Wgt_8_402,.Wgt_8_403,.Wgt_8_404,.Wgt_8_405,.Wgt_8_406,.Wgt_8_407,.Wgt_8_408,.Wgt_8_409,.Wgt_8_410,.Wgt_8_411,.Wgt_8_412,.Wgt_8_413,.Wgt_8_414,.Wgt_8_415,.Wgt_8_416,.Wgt_8_417,.Wgt_8_418,.Wgt_8_419,.Wgt_8_420,.Wgt_8_421,.Wgt_8_422,.Wgt_8_423,.Wgt_8_424,.Wgt_8_425,.Wgt_8_426,.Wgt_8_427,.Wgt_8_428,.Wgt_8_429,.Wgt_8_430,.Wgt_8_431,.Wgt_8_432,.Wgt_8_433,.Wgt_8_434,.Wgt_8_435,.Wgt_8_436,.Wgt_8_437,.Wgt_8_438,.Wgt_8_439,.Wgt_8_440,.Wgt_8_441,.Wgt_8_442,.Wgt_8_443,.Wgt_8_444,.Wgt_8_445,.Wgt_8_446,.Wgt_8_447,.Wgt_8_448,.Wgt_8_449,.Wgt_8_450,.Wgt_8_451,.Wgt_8_452,.Wgt_8_453,.Wgt_8_454,.Wgt_8_455,.Wgt_8_456,.Wgt_8_457,.Wgt_8_458,.Wgt_8_459,.Wgt_8_460,.Wgt_8_461,.Wgt_8_462,.Wgt_8_463,.Wgt_8_464,.Wgt_8_465,.Wgt_8_466,.Wgt_8_467,.Wgt_8_468,.Wgt_8_469,.Wgt_8_470,.Wgt_8_471,.Wgt_8_472,.Wgt_8_473,.Wgt_8_474,.Wgt_8_475,.Wgt_8_476,.Wgt_8_477,.Wgt_8_478,.Wgt_8_479,.Wgt_8_480,.Wgt_8_481,.Wgt_8_482,.Wgt_8_483,.Wgt_8_484,.Wgt_8_485,.Wgt_8_486,.Wgt_8_487,.Wgt_8_488,.Wgt_8_489,.Wgt_8_490,.Wgt_8_491,.Wgt_8_492,.Wgt_8_493,.Wgt_8_494,.Wgt_8_495,.Wgt_8_496,.Wgt_8_497,.Wgt_8_498,.Wgt_8_499,.Wgt_8_500,.Wgt_8_501,.Wgt_8_502,.Wgt_8_503,.Wgt_8_504,.Wgt_8_505,.Wgt_8_506,.Wgt_8_507,.Wgt_8_508,.Wgt_8_509,.Wgt_8_510,.Wgt_8_511,.Wgt_8_512,.Wgt_8_513,.Wgt_8_514,.Wgt_8_515,.Wgt_8_516,.Wgt_8_517,.Wgt_8_518,.Wgt_8_519,.Wgt_8_520,.Wgt_8_521,.Wgt_8_522,.Wgt_8_523,.Wgt_8_524,.Wgt_8_525,.Wgt_8_526,.Wgt_8_527,.Wgt_8_528,.Wgt_8_529,.Wgt_8_530,.Wgt_8_531,.Wgt_8_532,.Wgt_8_533,.Wgt_8_534,.Wgt_8_535,.Wgt_8_536,.Wgt_8_537,.Wgt_8_538,.Wgt_8_539,.Wgt_8_540,.Wgt_8_541,.Wgt_8_542,.Wgt_8_543,.Wgt_8_544,.Wgt_8_545,.Wgt_8_546,.Wgt_8_547,.Wgt_8_548,.Wgt_8_549,.Wgt_8_550,.Wgt_8_551,.Wgt_8_552,.Wgt_8_553,.Wgt_8_554,.Wgt_8_555,.Wgt_8_556,.Wgt_8_557,.Wgt_8_558,.Wgt_8_559,.Wgt_8_560,.Wgt_8_561,.Wgt_8_562,.Wgt_8_563,.Wgt_8_564,.Wgt_8_565,.Wgt_8_566,.Wgt_8_567,.Wgt_8_568,.Wgt_8_569,.Wgt_8_570,.Wgt_8_571,.Wgt_8_572,.Wgt_8_573,.Wgt_8_574,.Wgt_8_575,.Wgt_8_576,.Wgt_8_577,.Wgt_8_578,.Wgt_8_579,.Wgt_8_580,.Wgt_8_581,.Wgt_8_582,.Wgt_8_583,.Wgt_8_584,.Wgt_8_585,.Wgt_8_586,.Wgt_8_587,.Wgt_8_588,.Wgt_8_589,.Wgt_8_590,.Wgt_8_591,.Wgt_8_592,.Wgt_8_593,.Wgt_8_594,.Wgt_8_595,.Wgt_8_596,.Wgt_8_597,.Wgt_8_598,.Wgt_8_599,.Wgt_8_600,.Wgt_8_601,.Wgt_8_602,.Wgt_8_603,.Wgt_8_604,.Wgt_8_605,.Wgt_8_606,.Wgt_8_607,.Wgt_8_608,.Wgt_8_609,.Wgt_8_610,.Wgt_8_611,.Wgt_8_612,.Wgt_8_613,.Wgt_8_614,.Wgt_8_615,.Wgt_8_616,.Wgt_8_617,.Wgt_8_618,.Wgt_8_619,.Wgt_8_620,.Wgt_8_621,.Wgt_8_622,.Wgt_8_623,.Wgt_8_624,.Wgt_8_625,.Wgt_8_626,.Wgt_8_627,.Wgt_8_628,.Wgt_8_629,.Wgt_8_630,.Wgt_8_631,.Wgt_8_632,.Wgt_8_633,.Wgt_8_634,.Wgt_8_635,.Wgt_8_636,.Wgt_8_637,.Wgt_8_638,.Wgt_8_639,.Wgt_8_640,.Wgt_8_641,.Wgt_8_642,.Wgt_8_643,.Wgt_8_644,.Wgt_8_645,.Wgt_8_646,.Wgt_8_647,.Wgt_8_648,.Wgt_8_649,.Wgt_8_650,.Wgt_8_651,.Wgt_8_652,.Wgt_8_653,.Wgt_8_654,.Wgt_8_655,.Wgt_8_656,.Wgt_8_657,.Wgt_8_658,.Wgt_8_659,.Wgt_8_660,.Wgt_8_661,.Wgt_8_662,.Wgt_8_663,.Wgt_8_664,.Wgt_8_665,.Wgt_8_666,.Wgt_8_667,.Wgt_8_668,.Wgt_8_669,.Wgt_8_670,.Wgt_8_671,.Wgt_8_672,.Wgt_8_673,.Wgt_8_674,.Wgt_8_675,.Wgt_8_676,.Wgt_8_677,.Wgt_8_678,.Wgt_8_679,.Wgt_8_680,.Wgt_8_681,.Wgt_8_682,.Wgt_8_683,.Wgt_8_684,.Wgt_8_685,.Wgt_8_686,.Wgt_8_687,.Wgt_8_688,.Wgt_8_689,.Wgt_8_690,.Wgt_8_691,.Wgt_8_692,.Wgt_8_693,.Wgt_8_694,.Wgt_8_695,.Wgt_8_696,.Wgt_8_697,.Wgt_8_698,.Wgt_8_699,.Wgt_8_700,.Wgt_8_701,.Wgt_8_702,.Wgt_8_703,.Wgt_8_704,.Wgt_8_705,.Wgt_8_706,.Wgt_8_707,.Wgt_8_708,.Wgt_8_709,.Wgt_8_710,.Wgt_8_711,.Wgt_8_712,.Wgt_8_713,.Wgt_8_714,.Wgt_8_715,.Wgt_8_716,.Wgt_8_717,.Wgt_8_718,.Wgt_8_719,.Wgt_8_720,.Wgt_8_721,.Wgt_8_722,.Wgt_8_723,.Wgt_8_724,.Wgt_8_725,.Wgt_8_726,.Wgt_8_727,.Wgt_8_728,.Wgt_8_729,.Wgt_8_730,.Wgt_8_731,.Wgt_8_732,.Wgt_8_733,.Wgt_8_734,.Wgt_8_735,.Wgt_8_736,.Wgt_8_737,.Wgt_8_738,.Wgt_8_739,.Wgt_8_740,.Wgt_8_741,.Wgt_8_742,.Wgt_8_743,.Wgt_8_744,.Wgt_8_745,.Wgt_8_746,.Wgt_8_747,.Wgt_8_748,.Wgt_8_749,.Wgt_8_750,.Wgt_8_751,.Wgt_8_752,.Wgt_8_753,.Wgt_8_754,.Wgt_8_755,.Wgt_8_756,.Wgt_8_757,.Wgt_8_758,.Wgt_8_759,.Wgt_8_760,.Wgt_8_761,.Wgt_8_762,.Wgt_8_763,.Wgt_8_764,.Wgt_8_765,.Wgt_8_766,.Wgt_8_767,.Wgt_8_768,.Wgt_8_769,.Wgt_8_770,.Wgt_8_771,.Wgt_8_772,.Wgt_8_773,.Wgt_8_774,.Wgt_8_775,.Wgt_8_776,.Wgt_8_777,.Wgt_8_778,.Wgt_8_779,.Wgt_8_780,.Wgt_8_781,.Wgt_8_782,.Wgt_8_783,.Wgt_8_784,
.Wgt_9_0,.Wgt_9_1,.Wgt_9_2,.Wgt_9_3,.Wgt_9_4,.Wgt_9_5,.Wgt_9_6,.Wgt_9_7,.Wgt_9_8,.Wgt_9_9,.Wgt_9_10,.Wgt_9_11,.Wgt_9_12,.Wgt_9_13,.Wgt_9_14,.Wgt_9_15,.Wgt_9_16,.Wgt_9_17,.Wgt_9_18,.Wgt_9_19,.Wgt_9_20,.Wgt_9_21,.Wgt_9_22,.Wgt_9_23,.Wgt_9_24,.Wgt_9_25,.Wgt_9_26,.Wgt_9_27,.Wgt_9_28,.Wgt_9_29,.Wgt_9_30,.Wgt_9_31,.Wgt_9_32,.Wgt_9_33,.Wgt_9_34,.Wgt_9_35,.Wgt_9_36,.Wgt_9_37,.Wgt_9_38,.Wgt_9_39,.Wgt_9_40,.Wgt_9_41,.Wgt_9_42,.Wgt_9_43,.Wgt_9_44,.Wgt_9_45,.Wgt_9_46,.Wgt_9_47,.Wgt_9_48,.Wgt_9_49,.Wgt_9_50,.Wgt_9_51,.Wgt_9_52,.Wgt_9_53,.Wgt_9_54,.Wgt_9_55,.Wgt_9_56,.Wgt_9_57,.Wgt_9_58,.Wgt_9_59,.Wgt_9_60,.Wgt_9_61,.Wgt_9_62,.Wgt_9_63,.Wgt_9_64,.Wgt_9_65,.Wgt_9_66,.Wgt_9_67,.Wgt_9_68,.Wgt_9_69,.Wgt_9_70,.Wgt_9_71,.Wgt_9_72,.Wgt_9_73,.Wgt_9_74,.Wgt_9_75,.Wgt_9_76,.Wgt_9_77,.Wgt_9_78,.Wgt_9_79,.Wgt_9_80,.Wgt_9_81,.Wgt_9_82,.Wgt_9_83,.Wgt_9_84,.Wgt_9_85,.Wgt_9_86,.Wgt_9_87,.Wgt_9_88,.Wgt_9_89,.Wgt_9_90,.Wgt_9_91,.Wgt_9_92,.Wgt_9_93,.Wgt_9_94,.Wgt_9_95,.Wgt_9_96,.Wgt_9_97,.Wgt_9_98,.Wgt_9_99,.Wgt_9_100,.Wgt_9_101,.Wgt_9_102,.Wgt_9_103,.Wgt_9_104,.Wgt_9_105,.Wgt_9_106,.Wgt_9_107,.Wgt_9_108,.Wgt_9_109,.Wgt_9_110,.Wgt_9_111,.Wgt_9_112,.Wgt_9_113,.Wgt_9_114,.Wgt_9_115,.Wgt_9_116,.Wgt_9_117,.Wgt_9_118,.Wgt_9_119,.Wgt_9_120,.Wgt_9_121,.Wgt_9_122,.Wgt_9_123,.Wgt_9_124,.Wgt_9_125,.Wgt_9_126,.Wgt_9_127,.Wgt_9_128,.Wgt_9_129,.Wgt_9_130,.Wgt_9_131,.Wgt_9_132,.Wgt_9_133,.Wgt_9_134,.Wgt_9_135,.Wgt_9_136,.Wgt_9_137,.Wgt_9_138,.Wgt_9_139,.Wgt_9_140,.Wgt_9_141,.Wgt_9_142,.Wgt_9_143,.Wgt_9_144,.Wgt_9_145,.Wgt_9_146,.Wgt_9_147,.Wgt_9_148,.Wgt_9_149,.Wgt_9_150,.Wgt_9_151,.Wgt_9_152,.Wgt_9_153,.Wgt_9_154,.Wgt_9_155,.Wgt_9_156,.Wgt_9_157,.Wgt_9_158,.Wgt_9_159,.Wgt_9_160,.Wgt_9_161,.Wgt_9_162,.Wgt_9_163,.Wgt_9_164,.Wgt_9_165,.Wgt_9_166,.Wgt_9_167,.Wgt_9_168,.Wgt_9_169,.Wgt_9_170,.Wgt_9_171,.Wgt_9_172,.Wgt_9_173,.Wgt_9_174,.Wgt_9_175,.Wgt_9_176,.Wgt_9_177,.Wgt_9_178,.Wgt_9_179,.Wgt_9_180,.Wgt_9_181,.Wgt_9_182,.Wgt_9_183,.Wgt_9_184,.Wgt_9_185,.Wgt_9_186,.Wgt_9_187,.Wgt_9_188,.Wgt_9_189,.Wgt_9_190,.Wgt_9_191,.Wgt_9_192,.Wgt_9_193,.Wgt_9_194,.Wgt_9_195,.Wgt_9_196,.Wgt_9_197,.Wgt_9_198,.Wgt_9_199,.Wgt_9_200,.Wgt_9_201,.Wgt_9_202,.Wgt_9_203,.Wgt_9_204,.Wgt_9_205,.Wgt_9_206,.Wgt_9_207,.Wgt_9_208,.Wgt_9_209,.Wgt_9_210,.Wgt_9_211,.Wgt_9_212,.Wgt_9_213,.Wgt_9_214,.Wgt_9_215,.Wgt_9_216,.Wgt_9_217,.Wgt_9_218,.Wgt_9_219,.Wgt_9_220,.Wgt_9_221,.Wgt_9_222,.Wgt_9_223,.Wgt_9_224,.Wgt_9_225,.Wgt_9_226,.Wgt_9_227,.Wgt_9_228,.Wgt_9_229,.Wgt_9_230,.Wgt_9_231,.Wgt_9_232,.Wgt_9_233,.Wgt_9_234,.Wgt_9_235,.Wgt_9_236,.Wgt_9_237,.Wgt_9_238,.Wgt_9_239,.Wgt_9_240,.Wgt_9_241,.Wgt_9_242,.Wgt_9_243,.Wgt_9_244,.Wgt_9_245,.Wgt_9_246,.Wgt_9_247,.Wgt_9_248,.Wgt_9_249,.Wgt_9_250,.Wgt_9_251,.Wgt_9_252,.Wgt_9_253,.Wgt_9_254,.Wgt_9_255,.Wgt_9_256,.Wgt_9_257,.Wgt_9_258,.Wgt_9_259,.Wgt_9_260,.Wgt_9_261,.Wgt_9_262,.Wgt_9_263,.Wgt_9_264,.Wgt_9_265,.Wgt_9_266,.Wgt_9_267,.Wgt_9_268,.Wgt_9_269,.Wgt_9_270,.Wgt_9_271,.Wgt_9_272,.Wgt_9_273,.Wgt_9_274,.Wgt_9_275,.Wgt_9_276,.Wgt_9_277,.Wgt_9_278,.Wgt_9_279,.Wgt_9_280,.Wgt_9_281,.Wgt_9_282,.Wgt_9_283,.Wgt_9_284,.Wgt_9_285,.Wgt_9_286,.Wgt_9_287,.Wgt_9_288,.Wgt_9_289,.Wgt_9_290,.Wgt_9_291,.Wgt_9_292,.Wgt_9_293,.Wgt_9_294,.Wgt_9_295,.Wgt_9_296,.Wgt_9_297,.Wgt_9_298,.Wgt_9_299,.Wgt_9_300,.Wgt_9_301,.Wgt_9_302,.Wgt_9_303,.Wgt_9_304,.Wgt_9_305,.Wgt_9_306,.Wgt_9_307,.Wgt_9_308,.Wgt_9_309,.Wgt_9_310,.Wgt_9_311,.Wgt_9_312,.Wgt_9_313,.Wgt_9_314,.Wgt_9_315,.Wgt_9_316,.Wgt_9_317,.Wgt_9_318,.Wgt_9_319,.Wgt_9_320,.Wgt_9_321,.Wgt_9_322,.Wgt_9_323,.Wgt_9_324,.Wgt_9_325,.Wgt_9_326,.Wgt_9_327,.Wgt_9_328,.Wgt_9_329,.Wgt_9_330,.Wgt_9_331,.Wgt_9_332,.Wgt_9_333,.Wgt_9_334,.Wgt_9_335,.Wgt_9_336,.Wgt_9_337,.Wgt_9_338,.Wgt_9_339,.Wgt_9_340,.Wgt_9_341,.Wgt_9_342,.Wgt_9_343,.Wgt_9_344,.Wgt_9_345,.Wgt_9_346,.Wgt_9_347,.Wgt_9_348,.Wgt_9_349,.Wgt_9_350,.Wgt_9_351,.Wgt_9_352,.Wgt_9_353,.Wgt_9_354,.Wgt_9_355,.Wgt_9_356,.Wgt_9_357,.Wgt_9_358,.Wgt_9_359,.Wgt_9_360,.Wgt_9_361,.Wgt_9_362,.Wgt_9_363,.Wgt_9_364,.Wgt_9_365,.Wgt_9_366,.Wgt_9_367,.Wgt_9_368,.Wgt_9_369,.Wgt_9_370,.Wgt_9_371,.Wgt_9_372,.Wgt_9_373,.Wgt_9_374,.Wgt_9_375,.Wgt_9_376,.Wgt_9_377,.Wgt_9_378,.Wgt_9_379,.Wgt_9_380,.Wgt_9_381,.Wgt_9_382,.Wgt_9_383,.Wgt_9_384,.Wgt_9_385,.Wgt_9_386,.Wgt_9_387,.Wgt_9_388,.Wgt_9_389,.Wgt_9_390,.Wgt_9_391,.Wgt_9_392,.Wgt_9_393,.Wgt_9_394,.Wgt_9_395,.Wgt_9_396,.Wgt_9_397,.Wgt_9_398,.Wgt_9_399,.Wgt_9_400,.Wgt_9_401,.Wgt_9_402,.Wgt_9_403,.Wgt_9_404,.Wgt_9_405,.Wgt_9_406,.Wgt_9_407,.Wgt_9_408,.Wgt_9_409,.Wgt_9_410,.Wgt_9_411,.Wgt_9_412,.Wgt_9_413,.Wgt_9_414,.Wgt_9_415,.Wgt_9_416,.Wgt_9_417,.Wgt_9_418,.Wgt_9_419,.Wgt_9_420,.Wgt_9_421,.Wgt_9_422,.Wgt_9_423,.Wgt_9_424,.Wgt_9_425,.Wgt_9_426,.Wgt_9_427,.Wgt_9_428,.Wgt_9_429,.Wgt_9_430,.Wgt_9_431,.Wgt_9_432,.Wgt_9_433,.Wgt_9_434,.Wgt_9_435,.Wgt_9_436,.Wgt_9_437,.Wgt_9_438,.Wgt_9_439,.Wgt_9_440,.Wgt_9_441,.Wgt_9_442,.Wgt_9_443,.Wgt_9_444,.Wgt_9_445,.Wgt_9_446,.Wgt_9_447,.Wgt_9_448,.Wgt_9_449,.Wgt_9_450,.Wgt_9_451,.Wgt_9_452,.Wgt_9_453,.Wgt_9_454,.Wgt_9_455,.Wgt_9_456,.Wgt_9_457,.Wgt_9_458,.Wgt_9_459,.Wgt_9_460,.Wgt_9_461,.Wgt_9_462,.Wgt_9_463,.Wgt_9_464,.Wgt_9_465,.Wgt_9_466,.Wgt_9_467,.Wgt_9_468,.Wgt_9_469,.Wgt_9_470,.Wgt_9_471,.Wgt_9_472,.Wgt_9_473,.Wgt_9_474,.Wgt_9_475,.Wgt_9_476,.Wgt_9_477,.Wgt_9_478,.Wgt_9_479,.Wgt_9_480,.Wgt_9_481,.Wgt_9_482,.Wgt_9_483,.Wgt_9_484,.Wgt_9_485,.Wgt_9_486,.Wgt_9_487,.Wgt_9_488,.Wgt_9_489,.Wgt_9_490,.Wgt_9_491,.Wgt_9_492,.Wgt_9_493,.Wgt_9_494,.Wgt_9_495,.Wgt_9_496,.Wgt_9_497,.Wgt_9_498,.Wgt_9_499,.Wgt_9_500,.Wgt_9_501,.Wgt_9_502,.Wgt_9_503,.Wgt_9_504,.Wgt_9_505,.Wgt_9_506,.Wgt_9_507,.Wgt_9_508,.Wgt_9_509,.Wgt_9_510,.Wgt_9_511,.Wgt_9_512,.Wgt_9_513,.Wgt_9_514,.Wgt_9_515,.Wgt_9_516,.Wgt_9_517,.Wgt_9_518,.Wgt_9_519,.Wgt_9_520,.Wgt_9_521,.Wgt_9_522,.Wgt_9_523,.Wgt_9_524,.Wgt_9_525,.Wgt_9_526,.Wgt_9_527,.Wgt_9_528,.Wgt_9_529,.Wgt_9_530,.Wgt_9_531,.Wgt_9_532,.Wgt_9_533,.Wgt_9_534,.Wgt_9_535,.Wgt_9_536,.Wgt_9_537,.Wgt_9_538,.Wgt_9_539,.Wgt_9_540,.Wgt_9_541,.Wgt_9_542,.Wgt_9_543,.Wgt_9_544,.Wgt_9_545,.Wgt_9_546,.Wgt_9_547,.Wgt_9_548,.Wgt_9_549,.Wgt_9_550,.Wgt_9_551,.Wgt_9_552,.Wgt_9_553,.Wgt_9_554,.Wgt_9_555,.Wgt_9_556,.Wgt_9_557,.Wgt_9_558,.Wgt_9_559,.Wgt_9_560,.Wgt_9_561,.Wgt_9_562,.Wgt_9_563,.Wgt_9_564,.Wgt_9_565,.Wgt_9_566,.Wgt_9_567,.Wgt_9_568,.Wgt_9_569,.Wgt_9_570,.Wgt_9_571,.Wgt_9_572,.Wgt_9_573,.Wgt_9_574,.Wgt_9_575,.Wgt_9_576,.Wgt_9_577,.Wgt_9_578,.Wgt_9_579,.Wgt_9_580,.Wgt_9_581,.Wgt_9_582,.Wgt_9_583,.Wgt_9_584,.Wgt_9_585,.Wgt_9_586,.Wgt_9_587,.Wgt_9_588,.Wgt_9_589,.Wgt_9_590,.Wgt_9_591,.Wgt_9_592,.Wgt_9_593,.Wgt_9_594,.Wgt_9_595,.Wgt_9_596,.Wgt_9_597,.Wgt_9_598,.Wgt_9_599,.Wgt_9_600,.Wgt_9_601,.Wgt_9_602,.Wgt_9_603,.Wgt_9_604,.Wgt_9_605,.Wgt_9_606,.Wgt_9_607,.Wgt_9_608,.Wgt_9_609,.Wgt_9_610,.Wgt_9_611,.Wgt_9_612,.Wgt_9_613,.Wgt_9_614,.Wgt_9_615,.Wgt_9_616,.Wgt_9_617,.Wgt_9_618,.Wgt_9_619,.Wgt_9_620,.Wgt_9_621,.Wgt_9_622,.Wgt_9_623,.Wgt_9_624,.Wgt_9_625,.Wgt_9_626,.Wgt_9_627,.Wgt_9_628,.Wgt_9_629,.Wgt_9_630,.Wgt_9_631,.Wgt_9_632,.Wgt_9_633,.Wgt_9_634,.Wgt_9_635,.Wgt_9_636,.Wgt_9_637,.Wgt_9_638,.Wgt_9_639,.Wgt_9_640,.Wgt_9_641,.Wgt_9_642,.Wgt_9_643,.Wgt_9_644,.Wgt_9_645,.Wgt_9_646,.Wgt_9_647,.Wgt_9_648,.Wgt_9_649,.Wgt_9_650,.Wgt_9_651,.Wgt_9_652,.Wgt_9_653,.Wgt_9_654,.Wgt_9_655,.Wgt_9_656,.Wgt_9_657,.Wgt_9_658,.Wgt_9_659,.Wgt_9_660,.Wgt_9_661,.Wgt_9_662,.Wgt_9_663,.Wgt_9_664,.Wgt_9_665,.Wgt_9_666,.Wgt_9_667,.Wgt_9_668,.Wgt_9_669,.Wgt_9_670,.Wgt_9_671,.Wgt_9_672,.Wgt_9_673,.Wgt_9_674,.Wgt_9_675,.Wgt_9_676,.Wgt_9_677,.Wgt_9_678,.Wgt_9_679,.Wgt_9_680,.Wgt_9_681,.Wgt_9_682,.Wgt_9_683,.Wgt_9_684,.Wgt_9_685,.Wgt_9_686,.Wgt_9_687,.Wgt_9_688,.Wgt_9_689,.Wgt_9_690,.Wgt_9_691,.Wgt_9_692,.Wgt_9_693,.Wgt_9_694,.Wgt_9_695,.Wgt_9_696,.Wgt_9_697,.Wgt_9_698,.Wgt_9_699,.Wgt_9_700,.Wgt_9_701,.Wgt_9_702,.Wgt_9_703,.Wgt_9_704,.Wgt_9_705,.Wgt_9_706,.Wgt_9_707,.Wgt_9_708,.Wgt_9_709,.Wgt_9_710,.Wgt_9_711,.Wgt_9_712,.Wgt_9_713,.Wgt_9_714,.Wgt_9_715,.Wgt_9_716,.Wgt_9_717,.Wgt_9_718,.Wgt_9_719,.Wgt_9_720,.Wgt_9_721,.Wgt_9_722,.Wgt_9_723,.Wgt_9_724,.Wgt_9_725,.Wgt_9_726,.Wgt_9_727,.Wgt_9_728,.Wgt_9_729,.Wgt_9_730,.Wgt_9_731,.Wgt_9_732,.Wgt_9_733,.Wgt_9_734,.Wgt_9_735,.Wgt_9_736,.Wgt_9_737,.Wgt_9_738,.Wgt_9_739,.Wgt_9_740,.Wgt_9_741,.Wgt_9_742,.Wgt_9_743,.Wgt_9_744,.Wgt_9_745,.Wgt_9_746,.Wgt_9_747,.Wgt_9_748,.Wgt_9_749,.Wgt_9_750,.Wgt_9_751,.Wgt_9_752,.Wgt_9_753,.Wgt_9_754,.Wgt_9_755,.Wgt_9_756,.Wgt_9_757,.Wgt_9_758,.Wgt_9_759,.Wgt_9_760,.Wgt_9_761,.Wgt_9_762,.Wgt_9_763,.Wgt_9_764,.Wgt_9_765,.Wgt_9_766,.Wgt_9_767,.Wgt_9_768,.Wgt_9_769,.Wgt_9_770,.Wgt_9_771,.Wgt_9_772,.Wgt_9_773,.Wgt_9_774,.Wgt_9_775,.Wgt_9_776,.Wgt_9_777,.Wgt_9_778,.Wgt_9_779,.Wgt_9_780,.Wgt_9_781,.Wgt_9_782,.Wgt_9_783,.Wgt_9_784,
.neuron_0_mul_0_w, .neuron_0_mul_1_w, .neuron_0_mul_2_w, .neuron_0_mul_3_w, .neuron_0_mul_4_w, .neuron_0_mul_5_w, .neuron_0_mul_6_w, .neuron_0_mul_7_w, .neuron_0_mul_8_w, .neuron_0_mul_9_w, .neuron_0_mul_10_w, .neuron_0_mul_11_w, .neuron_0_mul_12_w, .neuron_0_mul_13_w, .neuron_0_mul_14_w, .neuron_0_mul_15_w, .neuron_0_mul_16_w, .neuron_0_mul_17_w, .neuron_0_mul_18_w, .neuron_0_mul_19_w, .neuron_0_mul_20_w, .neuron_0_mul_21_w, .neuron_0_mul_22_w, .neuron_0_mul_23_w, .neuron_0_mul_24_w, .neuron_0_mul_25_w, .neuron_0_mul_26_w, .neuron_0_mul_27_w,
.neuron_1_mul_0_w, .neuron_1_mul_1_w, .neuron_1_mul_2_w, .neuron_1_mul_3_w, .neuron_1_mul_4_w, .neuron_1_mul_5_w, .neuron_1_mul_6_w, .neuron_1_mul_7_w, .neuron_1_mul_8_w, .neuron_1_mul_9_w, .neuron_1_mul_10_w, .neuron_1_mul_11_w, .neuron_1_mul_12_w, .neuron_1_mul_13_w, .neuron_1_mul_14_w, .neuron_1_mul_15_w, .neuron_1_mul_16_w, .neuron_1_mul_17_w, .neuron_1_mul_18_w, .neuron_1_mul_19_w, .neuron_1_mul_20_w, .neuron_1_mul_21_w, .neuron_1_mul_22_w, .neuron_1_mul_23_w, .neuron_1_mul_24_w, .neuron_1_mul_25_w, .neuron_1_mul_26_w, .neuron_1_mul_27_w,
.neuron_2_mul_0_w, .neuron_2_mul_1_w, .neuron_2_mul_2_w, .neuron_2_mul_3_w, .neuron_2_mul_4_w, .neuron_2_mul_5_w, .neuron_2_mul_6_w, .neuron_2_mul_7_w, .neuron_2_mul_8_w, .neuron_2_mul_9_w, .neuron_2_mul_10_w, .neuron_2_mul_11_w, .neuron_2_mul_12_w, .neuron_2_mul_13_w, .neuron_2_mul_14_w, .neuron_2_mul_15_w, .neuron_2_mul_16_w, .neuron_2_mul_17_w, .neuron_2_mul_18_w, .neuron_2_mul_19_w, .neuron_2_mul_20_w, .neuron_2_mul_21_w, .neuron_2_mul_22_w, .neuron_2_mul_23_w, .neuron_2_mul_24_w, .neuron_2_mul_25_w, .neuron_2_mul_26_w, .neuron_2_mul_27_w,
.neuron_3_mul_0_w, .neuron_3_mul_1_w, .neuron_3_mul_2_w, .neuron_3_mul_3_w, .neuron_3_mul_4_w, .neuron_3_mul_5_w, .neuron_3_mul_6_w, .neuron_3_mul_7_w, .neuron_3_mul_8_w, .neuron_3_mul_9_w, .neuron_3_mul_10_w, .neuron_3_mul_11_w, .neuron_3_mul_12_w, .neuron_3_mul_13_w, .neuron_3_mul_14_w, .neuron_3_mul_15_w, .neuron_3_mul_16_w, .neuron_3_mul_17_w, .neuron_3_mul_18_w, .neuron_3_mul_19_w, .neuron_3_mul_20_w, .neuron_3_mul_21_w, .neuron_3_mul_22_w, .neuron_3_mul_23_w, .neuron_3_mul_24_w, .neuron_3_mul_25_w, .neuron_3_mul_26_w, .neuron_3_mul_27_w,
.neuron_4_mul_0_w, .neuron_4_mul_1_w, .neuron_4_mul_2_w, .neuron_4_mul_3_w, .neuron_4_mul_4_w, .neuron_4_mul_5_w, .neuron_4_mul_6_w, .neuron_4_mul_7_w, .neuron_4_mul_8_w, .neuron_4_mul_9_w, .neuron_4_mul_10_w, .neuron_4_mul_11_w, .neuron_4_mul_12_w, .neuron_4_mul_13_w, .neuron_4_mul_14_w, .neuron_4_mul_15_w, .neuron_4_mul_16_w, .neuron_4_mul_17_w, .neuron_4_mul_18_w, .neuron_4_mul_19_w, .neuron_4_mul_20_w, .neuron_4_mul_21_w, .neuron_4_mul_22_w, .neuron_4_mul_23_w, .neuron_4_mul_24_w, .neuron_4_mul_25_w, .neuron_4_mul_26_w, .neuron_4_mul_27_w,
.neuron_5_mul_0_w, .neuron_5_mul_1_w, .neuron_5_mul_2_w, .neuron_5_mul_3_w, .neuron_5_mul_4_w, .neuron_5_mul_5_w, .neuron_5_mul_6_w, .neuron_5_mul_7_w, .neuron_5_mul_8_w, .neuron_5_mul_9_w, .neuron_5_mul_10_w, .neuron_5_mul_11_w, .neuron_5_mul_12_w, .neuron_5_mul_13_w, .neuron_5_mul_14_w, .neuron_5_mul_15_w, .neuron_5_mul_16_w, .neuron_5_mul_17_w, .neuron_5_mul_18_w, .neuron_5_mul_19_w, .neuron_5_mul_20_w, .neuron_5_mul_21_w, .neuron_5_mul_22_w, .neuron_5_mul_23_w, .neuron_5_mul_24_w, .neuron_5_mul_25_w, .neuron_5_mul_26_w, .neuron_5_mul_27_w,
.neuron_6_mul_0_w, .neuron_6_mul_1_w, .neuron_6_mul_2_w, .neuron_6_mul_3_w, .neuron_6_mul_4_w, .neuron_6_mul_5_w, .neuron_6_mul_6_w, .neuron_6_mul_7_w, .neuron_6_mul_8_w, .neuron_6_mul_9_w, .neuron_6_mul_10_w, .neuron_6_mul_11_w, .neuron_6_mul_12_w, .neuron_6_mul_13_w, .neuron_6_mul_14_w, .neuron_6_mul_15_w, .neuron_6_mul_16_w, .neuron_6_mul_17_w, .neuron_6_mul_18_w, .neuron_6_mul_19_w, .neuron_6_mul_20_w, .neuron_6_mul_21_w, .neuron_6_mul_22_w, .neuron_6_mul_23_w, .neuron_6_mul_24_w, .neuron_6_mul_25_w, .neuron_6_mul_26_w, .neuron_6_mul_27_w,
.neuron_7_mul_0_w, .neuron_7_mul_1_w, .neuron_7_mul_2_w, .neuron_7_mul_3_w, .neuron_7_mul_4_w, .neuron_7_mul_5_w, .neuron_7_mul_6_w, .neuron_7_mul_7_w, .neuron_7_mul_8_w, .neuron_7_mul_9_w, .neuron_7_mul_10_w, .neuron_7_mul_11_w, .neuron_7_mul_12_w, .neuron_7_mul_13_w, .neuron_7_mul_14_w, .neuron_7_mul_15_w, .neuron_7_mul_16_w, .neuron_7_mul_17_w, .neuron_7_mul_18_w, .neuron_7_mul_19_w, .neuron_7_mul_20_w, .neuron_7_mul_21_w, .neuron_7_mul_22_w, .neuron_7_mul_23_w, .neuron_7_mul_24_w, .neuron_7_mul_25_w, .neuron_7_mul_26_w, .neuron_7_mul_27_w,
.neuron_8_mul_0_w, .neuron_8_mul_1_w, .neuron_8_mul_2_w, .neuron_8_mul_3_w, .neuron_8_mul_4_w, .neuron_8_mul_5_w, .neuron_8_mul_6_w, .neuron_8_mul_7_w, .neuron_8_mul_8_w, .neuron_8_mul_9_w, .neuron_8_mul_10_w, .neuron_8_mul_11_w, .neuron_8_mul_12_w, .neuron_8_mul_13_w, .neuron_8_mul_14_w, .neuron_8_mul_15_w, .neuron_8_mul_16_w, .neuron_8_mul_17_w, .neuron_8_mul_18_w, .neuron_8_mul_19_w, .neuron_8_mul_20_w, .neuron_8_mul_21_w, .neuron_8_mul_22_w, .neuron_8_mul_23_w, .neuron_8_mul_24_w, .neuron_8_mul_25_w, .neuron_8_mul_26_w, .neuron_8_mul_27_w,
.neuron_9_mul_0_w, .neuron_9_mul_1_w, .neuron_9_mul_2_w, .neuron_9_mul_3_w, .neuron_9_mul_4_w, .neuron_9_mul_5_w, .neuron_9_mul_6_w, .neuron_9_mul_7_w, .neuron_9_mul_8_w, .neuron_9_mul_9_w, .neuron_9_mul_10_w, .neuron_9_mul_11_w, .neuron_9_mul_12_w, .neuron_9_mul_13_w, .neuron_9_mul_14_w, .neuron_9_mul_15_w, .neuron_9_mul_16_w, .neuron_9_mul_17_w, .neuron_9_mul_18_w, .neuron_9_mul_19_w, .neuron_9_mul_20_w, .neuron_9_mul_21_w, .neuron_9_mul_22_w, .neuron_9_mul_23_w, .neuron_9_mul_24_w, .neuron_9_mul_25_w, .neuron_9_mul_26_w, .neuron_9_mul_27_w
);

// Adder constraints: First edition, less effective
// Use N to control adder for more efficient operation
// neuron_0, Level 1: Multipliers to Adders, 14 adders needed
assign neuron_0_add_0_p1 = neuron_0_mul_0_out;
assign neuron_0_add_0_p2 = neuron_0_mul_1_out;
assign neuron_0_add_1_p1 = neuron_0_mul_2_out;
assign neuron_0_add_1_p2 = neuron_0_mul_3_out;
assign neuron_0_add_2_p1 = neuron_0_mul_4_out;
assign neuron_0_add_2_p2 = neuron_0_mul_5_out;
assign neuron_0_add_3_p1 = neuron_0_mul_6_out;
assign neuron_0_add_3_p2 = neuron_0_mul_7_out;
assign neuron_0_add_4_p1 = neuron_0_mul_8_out;
assign neuron_0_add_4_p2 = neuron_0_mul_9_out;
assign neuron_0_add_5_p1 = neuron_0_mul_10_out;
assign neuron_0_add_5_p2 = neuron_0_mul_11_out;
assign neuron_0_add_6_p1 = neuron_0_mul_12_out;
assign neuron_0_add_6_p2 = neuron_0_mul_13_out;
assign neuron_0_add_7_p1 = neuron_0_mul_14_out;
assign neuron_0_add_7_p2 = neuron_0_mul_15_out;
assign neuron_0_add_8_p1 = neuron_0_mul_16_out;
assign neuron_0_add_8_p2 = neuron_0_mul_17_out;
assign neuron_0_add_9_p1 = neuron_0_mul_18_out;
assign neuron_0_add_9_p2 = neuron_0_mul_19_out;
assign neuron_0_add_10_p1 = neuron_0_mul_20_out;
assign neuron_0_add_10_p2 = neuron_0_mul_21_out;
assign neuron_0_add_11_p1 = neuron_0_mul_22_out;
assign neuron_0_add_11_p2 = neuron_0_mul_23_out;
assign neuron_0_add_12_p1 = neuron_0_mul_24_out;
assign neuron_0_add_12_p2 = neuron_0_mul_25_out;
assign neuron_0_add_13_p1 = neuron_0_mul_26_out;
assign neuron_0_add_13_p2 = neuron_0_mul_27_out;
// neuron_0, Level 2: 7 adders needed
assign neuron_0_add_14_p1 = neuron_0_add_0_out;
assign neuron_0_add_14_p2 = neuron_0_add_1_out;
assign neuron_0_add_15_p1 = neuron_0_add_2_out;
assign neuron_0_add_15_p2 = neuron_0_add_3_out;
assign neuron_0_add_16_p1 = neuron_0_add_4_out;
assign neuron_0_add_16_p2 = neuron_0_add_5_out;
assign neuron_0_add_17_p1 = neuron_0_add_6_out;
assign neuron_0_add_17_p2 = neuron_0_add_7_out;
assign neuron_0_add_18_p1 = neuron_0_add_8_out;
assign neuron_0_add_18_p2 = neuron_0_add_9_out;
assign neuron_0_add_19_p1 = neuron_0_add_10_out;
assign neuron_0_add_19_p2 = neuron_0_add_11_out;
assign neuron_0_add_20_p1 = neuron_0_add_12_out;
assign neuron_0_add_20_p2 = neuron_0_add_13_out;
// neuron_0, Level 3: 4 adders needed
assign neuron_0_add_21_p1 = neuron_0_add_14_out;
assign neuron_0_add_21_p2 = neuron_0_add_15_out;
assign neuron_0_add_22_p1 = neuron_0_add_16_out;
assign neuron_0_add_22_p2 = neuron_0_add_17_out;
assign neuron_0_add_23_p1 = neuron_0_add_18_out;
assign neuron_0_add_23_p2 = neuron_0_add_19_out;
assign neuron_0_add_24_p1 = neuron_0_add_20_out;
assign neuron_0_add_24_p2 = 0;  // Clearly this can be improved. Should be reconsidered after have a clearer understanding of timing
// neuron_0, Level 4: 2 adders needed
assign neuron_0_add_25_p1 = neuron_0_add_21_out;
assign neuron_0_add_25_p2 = neuron_0_add_22_out;
assign neuron_0_add_26_p1 = neuron_0_add_23_out;
assign neuron_0_add_26_p2 = neuron_0_add_24_out;
// neuron_0, Level 5: 1 adder needed
assign neuron_0_add_27_p1 = neuron_0_add_25_out;
assign neuron_0_add_27_p2 = neuron_0_add_26_out;
// neuron_0_add_27_out is the neuron final result of adding and multiplying

// neuron_1, Level 1: Multipliers to Adders, 14 adders needed
assign neuron_1_add_0_p1 = neuron_1_mul_0_out;
assign neuron_1_add_0_p2 = neuron_1_mul_1_out;
assign neuron_1_add_1_p1 = neuron_1_mul_2_out;
assign neuron_1_add_1_p2 = neuron_1_mul_3_out;
assign neuron_1_add_2_p1 = neuron_1_mul_4_out;
assign neuron_1_add_2_p2 = neuron_1_mul_5_out;
assign neuron_1_add_3_p1 = neuron_1_mul_6_out;
assign neuron_1_add_3_p2 = neuron_1_mul_7_out;
assign neuron_1_add_4_p1 = neuron_1_mul_8_out;
assign neuron_1_add_4_p2 = neuron_1_mul_9_out;
assign neuron_1_add_5_p1 = neuron_1_mul_10_out;
assign neuron_1_add_5_p2 = neuron_1_mul_11_out;
assign neuron_1_add_6_p1 = neuron_1_mul_12_out;
assign neuron_1_add_6_p2 = neuron_1_mul_13_out;
assign neuron_1_add_7_p1 = neuron_1_mul_14_out;
assign neuron_1_add_7_p2 = neuron_1_mul_15_out;
assign neuron_1_add_8_p1 = neuron_1_mul_16_out;
assign neuron_1_add_8_p2 = neuron_1_mul_17_out;
assign neuron_1_add_9_p1 = neuron_1_mul_18_out;
assign neuron_1_add_9_p2 = neuron_1_mul_19_out;
assign neuron_1_add_10_p1 = neuron_1_mul_20_out;
assign neuron_1_add_10_p2 = neuron_1_mul_21_out;
assign neuron_1_add_11_p1 = neuron_1_mul_22_out;
assign neuron_1_add_11_p2 = neuron_1_mul_23_out;
assign neuron_1_add_12_p1 = neuron_1_mul_24_out;
assign neuron_1_add_12_p2 = neuron_1_mul_25_out;
assign neuron_1_add_13_p1 = neuron_1_mul_26_out;
assign neuron_1_add_13_p2 = neuron_1_mul_27_out;
// neuron_1, Level 2: 7 adders needed
assign neuron_1_add_14_p1 = neuron_1_add_0_out;
assign neuron_1_add_14_p2 = neuron_1_add_1_out;
assign neuron_1_add_15_p1 = neuron_1_add_2_out;
assign neuron_1_add_15_p2 = neuron_1_add_3_out;
assign neuron_1_add_16_p1 = neuron_1_add_4_out;
assign neuron_1_add_16_p2 = neuron_1_add_5_out;
assign neuron_1_add_17_p1 = neuron_1_add_6_out;
assign neuron_1_add_17_p2 = neuron_1_add_7_out;
assign neuron_1_add_18_p1 = neuron_1_add_8_out;
assign neuron_1_add_18_p2 = neuron_1_add_9_out;
assign neuron_1_add_19_p1 = neuron_1_add_10_out;
assign neuron_1_add_19_p2 = neuron_1_add_11_out;
assign neuron_1_add_20_p1 = neuron_1_add_12_out;
assign neuron_1_add_20_p2 = neuron_1_add_13_out;
// neuron_1, Level 3: 4 adders needed
assign neuron_1_add_21_p1 = neuron_1_add_14_out;
assign neuron_1_add_21_p2 = neuron_1_add_15_out;
assign neuron_1_add_22_p1 = neuron_1_add_16_out;
assign neuron_1_add_22_p2 = neuron_1_add_17_out;
assign neuron_1_add_23_p1 = neuron_1_add_18_out;
assign neuron_1_add_23_p2 = neuron_1_add_19_out;
assign neuron_1_add_24_p1 = neuron_1_add_20_out;
assign neuron_1_add_24_p2 = 0;
// neuron_1, Level 4: 2 adders needed
assign neuron_1_add_25_p1 = neuron_1_add_21_out;
assign neuron_1_add_25_p2 = neuron_1_add_22_out;
assign neuron_1_add_26_p1 = neuron_1_add_23_out;
assign neuron_1_add_26_p2 = neuron_1_add_24_out;
// neuron_1, Level 5: 1 adder needed
assign neuron_1_add_27_p1 = neuron_1_add_25_out;
assign neuron_1_add_27_p2 = neuron_1_add_26_out;
// neuron_1_add_27_out is the neuron final result of adding and multiplying

// neuron_2, Level 1: Multipliers to Adders, 14 adders needed
assign neuron_2_add_0_p1 = neuron_2_mul_0_out;
assign neuron_2_add_0_p2 = neuron_2_mul_1_out;
assign neuron_2_add_1_p1 = neuron_2_mul_2_out;
assign neuron_2_add_1_p2 = neuron_2_mul_3_out;
assign neuron_2_add_2_p1 = neuron_2_mul_4_out;
assign neuron_2_add_2_p2 = neuron_2_mul_5_out;
assign neuron_2_add_3_p1 = neuron_2_mul_6_out;
assign neuron_2_add_3_p2 = neuron_2_mul_7_out;
assign neuron_2_add_4_p1 = neuron_2_mul_8_out;
assign neuron_2_add_4_p2 = neuron_2_mul_9_out;
assign neuron_2_add_5_p1 = neuron_2_mul_10_out;
assign neuron_2_add_5_p2 = neuron_2_mul_11_out;
assign neuron_2_add_6_p1 = neuron_2_mul_12_out;
assign neuron_2_add_6_p2 = neuron_2_mul_13_out;
assign neuron_2_add_7_p1 = neuron_2_mul_14_out;
assign neuron_2_add_7_p2 = neuron_2_mul_15_out;
assign neuron_2_add_8_p1 = neuron_2_mul_16_out;
assign neuron_2_add_8_p2 = neuron_2_mul_17_out;
assign neuron_2_add_9_p1 = neuron_2_mul_18_out;
assign neuron_2_add_9_p2 = neuron_2_mul_19_out;
assign neuron_2_add_10_p1 = neuron_2_mul_20_out;
assign neuron_2_add_10_p2 = neuron_2_mul_21_out;
assign neuron_2_add_11_p1 = neuron_2_mul_22_out;
assign neuron_2_add_11_p2 = neuron_2_mul_23_out;
assign neuron_2_add_12_p1 = neuron_2_mul_24_out;
assign neuron_2_add_12_p2 = neuron_2_mul_25_out;
assign neuron_2_add_13_p1 = neuron_2_mul_26_out;
assign neuron_2_add_13_p2 = neuron_2_mul_27_out;
// neuron_2, Level 2: 7 adders needed
assign neuron_2_add_14_p1 = neuron_2_add_0_out;
assign neuron_2_add_14_p2 = neuron_2_add_1_out;
assign neuron_2_add_15_p1 = neuron_2_add_2_out;
assign neuron_2_add_15_p2 = neuron_2_add_3_out;
assign neuron_2_add_16_p1 = neuron_2_add_4_out;
assign neuron_2_add_16_p2 = neuron_2_add_5_out;
assign neuron_2_add_17_p1 = neuron_2_add_6_out;
assign neuron_2_add_17_p2 = neuron_2_add_7_out;
assign neuron_2_add_18_p1 = neuron_2_add_8_out;
assign neuron_2_add_18_p2 = neuron_2_add_9_out;
assign neuron_2_add_19_p1 = neuron_2_add_10_out;
assign neuron_2_add_19_p2 = neuron_2_add_11_out;
assign neuron_2_add_20_p1 = neuron_2_add_12_out;
assign neuron_2_add_20_p2 = neuron_2_add_13_out;
// neuron_2, Level 3: 4 adders needed
assign neuron_2_add_21_p1 = neuron_2_add_14_out;
assign neuron_2_add_21_p2 = neuron_2_add_15_out;
assign neuron_2_add_22_p1 = neuron_2_add_16_out;
assign neuron_2_add_22_p2 = neuron_2_add_17_out;
assign neuron_2_add_23_p1 = neuron_2_add_18_out;
assign neuron_2_add_23_p2 = neuron_2_add_19_out;
assign neuron_2_add_24_p1 = neuron_2_add_20_out;
assign neuron_2_add_24_p2 = 0;
// neuron_2, Level 4: 2 adders needed
assign neuron_2_add_25_p1 = neuron_2_add_21_out;
assign neuron_2_add_25_p2 = neuron_2_add_22_out;
assign neuron_2_add_26_p1 = neuron_2_add_23_out;
assign neuron_2_add_26_p2 = neuron_2_add_24_out;
// neuron_2, Level 5: 1 adder needed
assign neuron_2_add_27_p1 = neuron_2_add_25_out;
assign neuron_2_add_27_p2 = neuron_2_add_26_out;
// neuron_2_add_27_out is the neuron final result of adding and multiplying

// neuron_3, Level 1: Multipliers to Adders, 14 adders needed
assign neuron_3_add_0_p1 = neuron_3_mul_0_out;
assign neuron_3_add_0_p2 = neuron_3_mul_1_out;
assign neuron_3_add_1_p1 = neuron_3_mul_2_out;
assign neuron_3_add_1_p2 = neuron_3_mul_3_out;
assign neuron_3_add_2_p1 = neuron_3_mul_4_out;
assign neuron_3_add_2_p2 = neuron_3_mul_5_out;
assign neuron_3_add_3_p1 = neuron_3_mul_6_out;
assign neuron_3_add_3_p2 = neuron_3_mul_7_out;
assign neuron_3_add_4_p1 = neuron_3_mul_8_out;
assign neuron_3_add_4_p2 = neuron_3_mul_9_out;
assign neuron_3_add_5_p1 = neuron_3_mul_10_out;
assign neuron_3_add_5_p2 = neuron_3_mul_11_out;
assign neuron_3_add_6_p1 = neuron_3_mul_12_out;
assign neuron_3_add_6_p2 = neuron_3_mul_13_out;
assign neuron_3_add_7_p1 = neuron_3_mul_14_out;
assign neuron_3_add_7_p2 = neuron_3_mul_15_out;
assign neuron_3_add_8_p1 = neuron_3_mul_16_out;
assign neuron_3_add_8_p2 = neuron_3_mul_17_out;
assign neuron_3_add_9_p1 = neuron_3_mul_18_out;
assign neuron_3_add_9_p2 = neuron_3_mul_19_out;
assign neuron_3_add_10_p1 = neuron_3_mul_20_out;
assign neuron_3_add_10_p2 = neuron_3_mul_21_out;
assign neuron_3_add_11_p1 = neuron_3_mul_22_out;
assign neuron_3_add_11_p2 = neuron_3_mul_23_out;
assign neuron_3_add_12_p1 = neuron_3_mul_24_out;
assign neuron_3_add_12_p2 = neuron_3_mul_25_out;
assign neuron_3_add_13_p1 = neuron_3_mul_26_out;
assign neuron_3_add_13_p2 = neuron_3_mul_27_out;
// neuron_3, Level 2: 7 adders needed
assign neuron_3_add_14_p1 = neuron_3_add_0_out;
assign neuron_3_add_14_p2 = neuron_3_add_1_out;
assign neuron_3_add_15_p1 = neuron_3_add_2_out;
assign neuron_3_add_15_p2 = neuron_3_add_3_out;
assign neuron_3_add_16_p1 = neuron_3_add_4_out;
assign neuron_3_add_16_p2 = neuron_3_add_5_out;
assign neuron_3_add_17_p1 = neuron_3_add_6_out;
assign neuron_3_add_17_p2 = neuron_3_add_7_out;
assign neuron_3_add_18_p1 = neuron_3_add_8_out;
assign neuron_3_add_18_p2 = neuron_3_add_9_out;
assign neuron_3_add_19_p1 = neuron_3_add_10_out;
assign neuron_3_add_19_p2 = neuron_3_add_11_out;
assign neuron_3_add_20_p1 = neuron_3_add_12_out;
assign neuron_3_add_20_p2 = neuron_3_add_13_out;
// neuron_3, Level 3: 4 adders needed
assign neuron_3_add_21_p1 = neuron_3_add_14_out;
assign neuron_3_add_21_p2 = neuron_3_add_15_out;
assign neuron_3_add_22_p1 = neuron_3_add_16_out;
assign neuron_3_add_22_p2 = neuron_3_add_17_out;
assign neuron_3_add_23_p1 = neuron_3_add_18_out;
assign neuron_3_add_23_p2 = neuron_3_add_19_out;
assign neuron_3_add_24_p1 = neuron_3_add_20_out;
assign neuron_3_add_24_p2 = 0;
// neuron_3, Level 4: 2 adders needed
assign neuron_3_add_25_p1 = neuron_3_add_21_out;
assign neuron_3_add_25_p2 = neuron_3_add_22_out;
assign neuron_3_add_26_p1 = neuron_3_add_23_out;
assign neuron_3_add_26_p2 = neuron_3_add_24_out;
// neuron_3, Level 5: 1 adder needed
assign neuron_3_add_27_p1 = neuron_3_add_25_out;
assign neuron_3_add_27_p2 = neuron_3_add_26_out;
// neuron_3_add_27_out is the neuron final result of adding and multiplying

// neuron_4, Level 1: Multipliers to Adders, 14 adders needed
assign neuron_4_add_0_p1 = neuron_4_mul_0_out;
assign neuron_4_add_0_p2 = neuron_4_mul_1_out;
assign neuron_4_add_1_p1 = neuron_4_mul_2_out;
assign neuron_4_add_1_p2 = neuron_4_mul_3_out;
assign neuron_4_add_2_p1 = neuron_4_mul_4_out;
assign neuron_4_add_2_p2 = neuron_4_mul_5_out;
assign neuron_4_add_3_p1 = neuron_4_mul_6_out;
assign neuron_4_add_3_p2 = neuron_4_mul_7_out;
assign neuron_4_add_4_p1 = neuron_4_mul_8_out;
assign neuron_4_add_4_p2 = neuron_4_mul_9_out;
assign neuron_4_add_5_p1 = neuron_4_mul_10_out;
assign neuron_4_add_5_p2 = neuron_4_mul_11_out;
assign neuron_4_add_6_p1 = neuron_4_mul_12_out;
assign neuron_4_add_6_p2 = neuron_4_mul_13_out;
assign neuron_4_add_7_p1 = neuron_4_mul_14_out;
assign neuron_4_add_7_p2 = neuron_4_mul_15_out;
assign neuron_4_add_8_p1 = neuron_4_mul_16_out;
assign neuron_4_add_8_p2 = neuron_4_mul_17_out;
assign neuron_4_add_9_p1 = neuron_4_mul_18_out;
assign neuron_4_add_9_p2 = neuron_4_mul_19_out;
assign neuron_4_add_10_p1 = neuron_4_mul_20_out;
assign neuron_4_add_10_p2 = neuron_4_mul_21_out;
assign neuron_4_add_11_p1 = neuron_4_mul_22_out;
assign neuron_4_add_11_p2 = neuron_4_mul_23_out;
assign neuron_4_add_12_p1 = neuron_4_mul_24_out;
assign neuron_4_add_12_p2 = neuron_4_mul_25_out;
assign neuron_4_add_13_p1 = neuron_4_mul_26_out;
assign neuron_4_add_13_p2 = neuron_4_mul_27_out;
// neuron_4, Level 2: 7 adders needed
assign neuron_4_add_14_p1 = neuron_4_add_0_out;
assign neuron_4_add_14_p2 = neuron_4_add_1_out;
assign neuron_4_add_15_p1 = neuron_4_add_2_out;
assign neuron_4_add_15_p2 = neuron_4_add_3_out;
assign neuron_4_add_16_p1 = neuron_4_add_4_out;
assign neuron_4_add_16_p2 = neuron_4_add_5_out;
assign neuron_4_add_17_p1 = neuron_4_add_6_out;
assign neuron_4_add_17_p2 = neuron_4_add_7_out;
assign neuron_4_add_18_p1 = neuron_4_add_8_out;
assign neuron_4_add_18_p2 = neuron_4_add_9_out;
assign neuron_4_add_19_p1 = neuron_4_add_10_out;
assign neuron_4_add_19_p2 = neuron_4_add_11_out;
assign neuron_4_add_20_p1 = neuron_4_add_12_out;
assign neuron_4_add_20_p2 = neuron_4_add_13_out;
// neuron_4, Level 3: 4 adders needed
assign neuron_4_add_21_p1 = neuron_4_add_14_out;
assign neuron_4_add_21_p2 = neuron_4_add_15_out;
assign neuron_4_add_22_p1 = neuron_4_add_16_out;
assign neuron_4_add_22_p2 = neuron_4_add_17_out;
assign neuron_4_add_23_p1 = neuron_4_add_18_out;
assign neuron_4_add_23_p2 = neuron_4_add_19_out;
assign neuron_4_add_24_p1 = neuron_4_add_20_out;
assign neuron_4_add_24_p2 = 0;
// neuron_4, Level 4: 2 adders needed
assign neuron_4_add_25_p1 = neuron_4_add_21_out;
assign neuron_4_add_25_p2 = neuron_4_add_22_out;
assign neuron_4_add_26_p1 = neuron_4_add_23_out;
assign neuron_4_add_26_p2 = neuron_4_add_24_out;
// neuron_4, Level 5: 1 adder needed
assign neuron_4_add_27_p1 = neuron_4_add_25_out;
assign neuron_4_add_27_p2 = neuron_4_add_26_out;
// neuron_4_add_27_out is the neuron final result of adding and multiplying

// neuron_5, Level 1: Multipliers to Adders, 14 adders needed
assign neuron_5_add_0_p1 = neuron_5_mul_0_out;
assign neuron_5_add_0_p2 = neuron_5_mul_1_out;
assign neuron_5_add_1_p1 = neuron_5_mul_2_out;
assign neuron_5_add_1_p2 = neuron_5_mul_3_out;
assign neuron_5_add_2_p1 = neuron_5_mul_4_out;
assign neuron_5_add_2_p2 = neuron_5_mul_5_out;
assign neuron_5_add_3_p1 = neuron_5_mul_6_out;
assign neuron_5_add_3_p2 = neuron_5_mul_7_out;
assign neuron_5_add_4_p1 = neuron_5_mul_8_out;
assign neuron_5_add_4_p2 = neuron_5_mul_9_out;
assign neuron_5_add_5_p1 = neuron_5_mul_10_out;
assign neuron_5_add_5_p2 = neuron_5_mul_11_out;
assign neuron_5_add_6_p1 = neuron_5_mul_12_out;
assign neuron_5_add_6_p2 = neuron_5_mul_13_out;
assign neuron_5_add_7_p1 = neuron_5_mul_14_out;
assign neuron_5_add_7_p2 = neuron_5_mul_15_out;
assign neuron_5_add_8_p1 = neuron_5_mul_16_out;
assign neuron_5_add_8_p2 = neuron_5_mul_17_out;
assign neuron_5_add_9_p1 = neuron_5_mul_18_out;
assign neuron_5_add_9_p2 = neuron_5_mul_19_out;
assign neuron_5_add_10_p1 = neuron_5_mul_20_out;
assign neuron_5_add_10_p2 = neuron_5_mul_21_out;
assign neuron_5_add_11_p1 = neuron_5_mul_22_out;
assign neuron_5_add_11_p2 = neuron_5_mul_23_out;
assign neuron_5_add_12_p1 = neuron_5_mul_24_out;
assign neuron_5_add_12_p2 = neuron_5_mul_25_out;
assign neuron_5_add_13_p1 = neuron_5_mul_26_out;
assign neuron_5_add_13_p2 = neuron_5_mul_27_out;
// neuron_5, Level 2: 7 adders needed
assign neuron_5_add_14_p1 = neuron_5_add_0_out;
assign neuron_5_add_14_p2 = neuron_5_add_1_out;
assign neuron_5_add_15_p1 = neuron_5_add_2_out;
assign neuron_5_add_15_p2 = neuron_5_add_3_out;
assign neuron_5_add_16_p1 = neuron_5_add_4_out;
assign neuron_5_add_16_p2 = neuron_5_add_5_out;
assign neuron_5_add_17_p1 = neuron_5_add_6_out;
assign neuron_5_add_17_p2 = neuron_5_add_7_out;
assign neuron_5_add_18_p1 = neuron_5_add_8_out;
assign neuron_5_add_18_p2 = neuron_5_add_9_out;
assign neuron_5_add_19_p1 = neuron_5_add_10_out;
assign neuron_5_add_19_p2 = neuron_5_add_11_out;
assign neuron_5_add_20_p1 = neuron_5_add_12_out;
assign neuron_5_add_20_p2 = neuron_5_add_13_out;
// neuron_5, Level 3: 4 adders needed
assign neuron_5_add_21_p1 = neuron_5_add_14_out;
assign neuron_5_add_21_p2 = neuron_5_add_15_out;
assign neuron_5_add_22_p1 = neuron_5_add_16_out;
assign neuron_5_add_22_p2 = neuron_5_add_17_out;
assign neuron_5_add_23_p1 = neuron_5_add_18_out;
assign neuron_5_add_23_p2 = neuron_5_add_19_out;
assign neuron_5_add_24_p1 = neuron_5_add_20_out;
assign neuron_5_add_24_p2 = 0;
// neuron_5, Level 4: 2 adders needed
assign neuron_5_add_25_p1 = neuron_5_add_21_out;
assign neuron_5_add_25_p2 = neuron_5_add_22_out;
assign neuron_5_add_26_p1 = neuron_5_add_23_out;
assign neuron_5_add_26_p2 = neuron_5_add_24_out;
// neuron_5, Level 5: 1 adder needed
assign neuron_5_add_27_p1 = neuron_5_add_25_out;
assign neuron_5_add_27_p2 = neuron_5_add_26_out;
// neuron_5_add_27_out is the neuron final result of adding and multiplying

// neuron_6, Level 1: Multipliers to Adders, 14 adders needed
assign neuron_6_add_0_p1 = neuron_6_mul_0_out;
assign neuron_6_add_0_p2 = neuron_6_mul_1_out;
assign neuron_6_add_1_p1 = neuron_6_mul_2_out;
assign neuron_6_add_1_p2 = neuron_6_mul_3_out;
assign neuron_6_add_2_p1 = neuron_6_mul_4_out;
assign neuron_6_add_2_p2 = neuron_6_mul_5_out;
assign neuron_6_add_3_p1 = neuron_6_mul_6_out;
assign neuron_6_add_3_p2 = neuron_6_mul_7_out;
assign neuron_6_add_4_p1 = neuron_6_mul_8_out;
assign neuron_6_add_4_p2 = neuron_6_mul_9_out;
assign neuron_6_add_5_p1 = neuron_6_mul_10_out;
assign neuron_6_add_5_p2 = neuron_6_mul_11_out;
assign neuron_6_add_6_p1 = neuron_6_mul_12_out;
assign neuron_6_add_6_p2 = neuron_6_mul_13_out;
assign neuron_6_add_7_p1 = neuron_6_mul_14_out;
assign neuron_6_add_7_p2 = neuron_6_mul_15_out;
assign neuron_6_add_8_p1 = neuron_6_mul_16_out;
assign neuron_6_add_8_p2 = neuron_6_mul_17_out;
assign neuron_6_add_9_p1 = neuron_6_mul_18_out;
assign neuron_6_add_9_p2 = neuron_6_mul_19_out;
assign neuron_6_add_10_p1 = neuron_6_mul_20_out;
assign neuron_6_add_10_p2 = neuron_6_mul_21_out;
assign neuron_6_add_11_p1 = neuron_6_mul_22_out;
assign neuron_6_add_11_p2 = neuron_6_mul_23_out;
assign neuron_6_add_12_p1 = neuron_6_mul_24_out;
assign neuron_6_add_12_p2 = neuron_6_mul_25_out;
assign neuron_6_add_13_p1 = neuron_6_mul_26_out;
assign neuron_6_add_13_p2 = neuron_6_mul_27_out;
// neuron_6, Level 2: 7 adders needed
assign neuron_6_add_14_p1 = neuron_6_add_0_out;
assign neuron_6_add_14_p2 = neuron_6_add_1_out;
assign neuron_6_add_15_p1 = neuron_6_add_2_out;
assign neuron_6_add_15_p2 = neuron_6_add_3_out;
assign neuron_6_add_16_p1 = neuron_6_add_4_out;
assign neuron_6_add_16_p2 = neuron_6_add_5_out;
assign neuron_6_add_17_p1 = neuron_6_add_6_out;
assign neuron_6_add_17_p2 = neuron_6_add_7_out;
assign neuron_6_add_18_p1 = neuron_6_add_8_out;
assign neuron_6_add_18_p2 = neuron_6_add_9_out;
assign neuron_6_add_19_p1 = neuron_6_add_10_out;
assign neuron_6_add_19_p2 = neuron_6_add_11_out;
assign neuron_6_add_20_p1 = neuron_6_add_12_out;
assign neuron_6_add_20_p2 = neuron_6_add_13_out;
// neuron_6, Level 3: 4 adders needed
assign neuron_6_add_21_p1 = neuron_6_add_14_out;
assign neuron_6_add_21_p2 = neuron_6_add_15_out;
assign neuron_6_add_22_p1 = neuron_6_add_16_out;
assign neuron_6_add_22_p2 = neuron_6_add_17_out;
assign neuron_6_add_23_p1 = neuron_6_add_18_out;
assign neuron_6_add_23_p2 = neuron_6_add_19_out;
assign neuron_6_add_24_p1 = neuron_6_add_20_out;
assign neuron_6_add_24_p2 = 0;
// neuron_6, Level 4: 2 adders needed
assign neuron_6_add_25_p1 = neuron_6_add_21_out;
assign neuron_6_add_25_p2 = neuron_6_add_22_out;
assign neuron_6_add_26_p1 = neuron_6_add_23_out;
assign neuron_6_add_26_p2 = neuron_6_add_24_out;
// neuron_6, Level 5: 1 adder needed
assign neuron_6_add_27_p1 = neuron_6_add_25_out;
assign neuron_6_add_27_p2 = neuron_6_add_26_out;
// neuron_6_add_27_out is the neuron final result of adding and multiplying

// neuron_7, Level 1: Multipliers to Adders, 14 adders needed
assign neuron_7_add_0_p1 = neuron_7_mul_0_out;
assign neuron_7_add_0_p2 = neuron_7_mul_1_out;
assign neuron_7_add_1_p1 = neuron_7_mul_2_out;
assign neuron_7_add_1_p2 = neuron_7_mul_3_out;
assign neuron_7_add_2_p1 = neuron_7_mul_4_out;
assign neuron_7_add_2_p2 = neuron_7_mul_5_out;
assign neuron_7_add_3_p1 = neuron_7_mul_6_out;
assign neuron_7_add_3_p2 = neuron_7_mul_7_out;
assign neuron_7_add_4_p1 = neuron_7_mul_8_out;
assign neuron_7_add_4_p2 = neuron_7_mul_9_out;
assign neuron_7_add_5_p1 = neuron_7_mul_10_out;
assign neuron_7_add_5_p2 = neuron_7_mul_11_out;
assign neuron_7_add_6_p1 = neuron_7_mul_12_out;
assign neuron_7_add_6_p2 = neuron_7_mul_13_out;
assign neuron_7_add_7_p1 = neuron_7_mul_14_out;
assign neuron_7_add_7_p2 = neuron_7_mul_15_out;
assign neuron_7_add_8_p1 = neuron_7_mul_16_out;
assign neuron_7_add_8_p2 = neuron_7_mul_17_out;
assign neuron_7_add_9_p1 = neuron_7_mul_18_out;
assign neuron_7_add_9_p2 = neuron_7_mul_19_out;
assign neuron_7_add_10_p1 = neuron_7_mul_20_out;
assign neuron_7_add_10_p2 = neuron_7_mul_21_out;
assign neuron_7_add_11_p1 = neuron_7_mul_22_out;
assign neuron_7_add_11_p2 = neuron_7_mul_23_out;
assign neuron_7_add_12_p1 = neuron_7_mul_24_out;
assign neuron_7_add_12_p2 = neuron_7_mul_25_out;
assign neuron_7_add_13_p1 = neuron_7_mul_26_out;
assign neuron_7_add_13_p2 = neuron_7_mul_27_out;
// neuron_7, Level 2: 7 adders needed
assign neuron_7_add_14_p1 = neuron_7_add_0_out;
assign neuron_7_add_14_p2 = neuron_7_add_1_out;
assign neuron_7_add_15_p1 = neuron_7_add_2_out;
assign neuron_7_add_15_p2 = neuron_7_add_3_out;
assign neuron_7_add_16_p1 = neuron_7_add_4_out;
assign neuron_7_add_16_p2 = neuron_7_add_5_out;
assign neuron_7_add_17_p1 = neuron_7_add_6_out;
assign neuron_7_add_17_p2 = neuron_7_add_7_out;
assign neuron_7_add_18_p1 = neuron_7_add_8_out;
assign neuron_7_add_18_p2 = neuron_7_add_9_out;
assign neuron_7_add_19_p1 = neuron_7_add_10_out;
assign neuron_7_add_19_p2 = neuron_7_add_11_out;
assign neuron_7_add_20_p1 = neuron_7_add_12_out;
assign neuron_7_add_20_p2 = neuron_7_add_13_out;
// neuron_7, Level 3: 4 adders needed
assign neuron_7_add_21_p1 = neuron_7_add_14_out;
assign neuron_7_add_21_p2 = neuron_7_add_15_out;
assign neuron_7_add_22_p1 = neuron_7_add_16_out;
assign neuron_7_add_22_p2 = neuron_7_add_17_out;
assign neuron_7_add_23_p1 = neuron_7_add_18_out;
assign neuron_7_add_23_p2 = neuron_7_add_19_out;
assign neuron_7_add_24_p1 = neuron_7_add_20_out;
assign neuron_7_add_24_p2 = 0;
// neuron_7, Level 4: 2 adders needed
assign neuron_7_add_25_p1 = neuron_7_add_21_out;
assign neuron_7_add_25_p2 = neuron_7_add_22_out;
assign neuron_7_add_26_p1 = neuron_7_add_23_out;
assign neuron_7_add_26_p2 = neuron_7_add_24_out;
// neuron_7, Level 5: 1 adder needed
assign neuron_7_add_27_p1 = neuron_7_add_25_out;
assign neuron_7_add_27_p2 = neuron_7_add_26_out;
// neuron_7_add_27_out is the neuron final result of adding and multiplying

// neuron_8, Level 1: Multipliers to Adders, 14 adders needed
assign neuron_8_add_0_p1 = neuron_8_mul_0_out;
assign neuron_8_add_0_p2 = neuron_8_mul_1_out;
assign neuron_8_add_1_p1 = neuron_8_mul_2_out;
assign neuron_8_add_1_p2 = neuron_8_mul_3_out;
assign neuron_8_add_2_p1 = neuron_8_mul_4_out;
assign neuron_8_add_2_p2 = neuron_8_mul_5_out;
assign neuron_8_add_3_p1 = neuron_8_mul_6_out;
assign neuron_8_add_3_p2 = neuron_8_mul_7_out;
assign neuron_8_add_4_p1 = neuron_8_mul_8_out;
assign neuron_8_add_4_p2 = neuron_8_mul_9_out;
assign neuron_8_add_5_p1 = neuron_8_mul_10_out;
assign neuron_8_add_5_p2 = neuron_8_mul_11_out;
assign neuron_8_add_6_p1 = neuron_8_mul_12_out;
assign neuron_8_add_6_p2 = neuron_8_mul_13_out;
assign neuron_8_add_7_p1 = neuron_8_mul_14_out;
assign neuron_8_add_7_p2 = neuron_8_mul_15_out;
assign neuron_8_add_8_p1 = neuron_8_mul_16_out;
assign neuron_8_add_8_p2 = neuron_8_mul_17_out;
assign neuron_8_add_9_p1 = neuron_8_mul_18_out;
assign neuron_8_add_9_p2 = neuron_8_mul_19_out;
assign neuron_8_add_10_p1 = neuron_8_mul_20_out;
assign neuron_8_add_10_p2 = neuron_8_mul_21_out;
assign neuron_8_add_11_p1 = neuron_8_mul_22_out;
assign neuron_8_add_11_p2 = neuron_8_mul_23_out;
assign neuron_8_add_12_p1 = neuron_8_mul_24_out;
assign neuron_8_add_12_p2 = neuron_8_mul_25_out;
assign neuron_8_add_13_p1 = neuron_8_mul_26_out;
assign neuron_8_add_13_p2 = neuron_8_mul_27_out;
// neuron_8, Level 2: 7 adders needed
assign neuron_8_add_14_p1 = neuron_8_add_0_out;
assign neuron_8_add_14_p2 = neuron_8_add_1_out;
assign neuron_8_add_15_p1 = neuron_8_add_2_out;
assign neuron_8_add_15_p2 = neuron_8_add_3_out;
assign neuron_8_add_16_p1 = neuron_8_add_4_out;
assign neuron_8_add_16_p2 = neuron_8_add_5_out;
assign neuron_8_add_17_p1 = neuron_8_add_6_out;
assign neuron_8_add_17_p2 = neuron_8_add_7_out;
assign neuron_8_add_18_p1 = neuron_8_add_8_out;
assign neuron_8_add_18_p2 = neuron_8_add_9_out;
assign neuron_8_add_19_p1 = neuron_8_add_10_out;
assign neuron_8_add_19_p2 = neuron_8_add_11_out;
assign neuron_8_add_20_p1 = neuron_8_add_12_out;
assign neuron_8_add_20_p2 = neuron_8_add_13_out;
// neuron_8, Level 3: 4 adders needed
assign neuron_8_add_21_p1 = neuron_8_add_14_out;
assign neuron_8_add_21_p2 = neuron_8_add_15_out;
assign neuron_8_add_22_p1 = neuron_8_add_16_out;
assign neuron_8_add_22_p2 = neuron_8_add_17_out;
assign neuron_8_add_23_p1 = neuron_8_add_18_out;
assign neuron_8_add_23_p2 = neuron_8_add_19_out;
assign neuron_8_add_24_p1 = neuron_8_add_20_out;
assign neuron_8_add_24_p2 = 0;
// neuron_8, Level 4: 2 adders needed
assign neuron_8_add_25_p1 = neuron_8_add_21_out;
assign neuron_8_add_25_p2 = neuron_8_add_22_out;
assign neuron_8_add_26_p1 = neuron_8_add_23_out;
assign neuron_8_add_26_p2 = neuron_8_add_24_out;
// neuron_8, Level 5: 1 adder needed
assign neuron_8_add_27_p1 = neuron_8_add_25_out;
assign neuron_8_add_27_p2 = neuron_8_add_26_out;
// neuron_8_add_27_out is the neuron final result of adding and multiplying

// neuron_9, Level 1: Multipliers to Adders, 14 adders needed
assign neuron_9_add_0_p1 = neuron_9_mul_0_out;
assign neuron_9_add_0_p2 = neuron_9_mul_1_out;
assign neuron_9_add_1_p1 = neuron_9_mul_2_out;
assign neuron_9_add_1_p2 = neuron_9_mul_3_out;
assign neuron_9_add_2_p1 = neuron_9_mul_4_out;
assign neuron_9_add_2_p2 = neuron_9_mul_5_out;
assign neuron_9_add_3_p1 = neuron_9_mul_6_out;
assign neuron_9_add_3_p2 = neuron_9_mul_7_out;
assign neuron_9_add_4_p1 = neuron_9_mul_8_out;
assign neuron_9_add_4_p2 = neuron_9_mul_9_out;
assign neuron_9_add_5_p1 = neuron_9_mul_10_out;
assign neuron_9_add_5_p2 = neuron_9_mul_11_out;
assign neuron_9_add_6_p1 = neuron_9_mul_12_out;
assign neuron_9_add_6_p2 = neuron_9_mul_13_out;
assign neuron_9_add_7_p1 = neuron_9_mul_14_out;
assign neuron_9_add_7_p2 = neuron_9_mul_15_out;
assign neuron_9_add_8_p1 = neuron_9_mul_16_out;
assign neuron_9_add_8_p2 = neuron_9_mul_17_out;
assign neuron_9_add_9_p1 = neuron_9_mul_18_out;
assign neuron_9_add_9_p2 = neuron_9_mul_19_out;
assign neuron_9_add_10_p1 = neuron_9_mul_20_out;
assign neuron_9_add_10_p2 = neuron_9_mul_21_out;
assign neuron_9_add_11_p1 = neuron_9_mul_22_out;
assign neuron_9_add_11_p2 = neuron_9_mul_23_out;
assign neuron_9_add_12_p1 = neuron_9_mul_24_out;
assign neuron_9_add_12_p2 = neuron_9_mul_25_out;
assign neuron_9_add_13_p1 = neuron_9_mul_26_out;
assign neuron_9_add_13_p2 = neuron_9_mul_27_out;
// neuron_9, Level 2: 7 adders needed
assign neuron_9_add_14_p1 = neuron_9_add_0_out;
assign neuron_9_add_14_p2 = neuron_9_add_1_out;
assign neuron_9_add_15_p1 = neuron_9_add_2_out;
assign neuron_9_add_15_p2 = neuron_9_add_3_out;
assign neuron_9_add_16_p1 = neuron_9_add_4_out;
assign neuron_9_add_16_p2 = neuron_9_add_5_out;
assign neuron_9_add_17_p1 = neuron_9_add_6_out;
assign neuron_9_add_17_p2 = neuron_9_add_7_out;
assign neuron_9_add_18_p1 = neuron_9_add_8_out;
assign neuron_9_add_18_p2 = neuron_9_add_9_out;
assign neuron_9_add_19_p1 = neuron_9_add_10_out;
assign neuron_9_add_19_p2 = neuron_9_add_11_out;
assign neuron_9_add_20_p1 = neuron_9_add_12_out;
assign neuron_9_add_20_p2 = neuron_9_add_13_out;
// neuron_9, Level 3: 4 adders needed
assign neuron_9_add_21_p1 = neuron_9_add_14_out;
assign neuron_9_add_21_p2 = neuron_9_add_15_out;
assign neuron_9_add_22_p1 = neuron_9_add_16_out;
assign neuron_9_add_22_p2 = neuron_9_add_17_out;
assign neuron_9_add_23_p1 = neuron_9_add_18_out;
assign neuron_9_add_23_p2 = neuron_9_add_19_out;
assign neuron_9_add_24_p1 = neuron_9_add_20_out;
assign neuron_9_add_24_p2 = 0;
// neuron_9, Level 4: 2 adders needed
assign neuron_9_add_25_p1 = neuron_9_add_21_out;
assign neuron_9_add_25_p2 = neuron_9_add_22_out;
assign neuron_9_add_26_p1 = neuron_9_add_23_out;
assign neuron_9_add_26_p2 = neuron_9_add_24_out;
// neuron_9, Level 5: 1 adder needed
assign neuron_9_add_27_p1 = neuron_9_add_25_out;
assign neuron_9_add_27_p2 = neuron_9_add_26_out;
// neuron_9_add_27_out is the neuron final result of adding and multiplying

// Final output of ten neurons
reg [25:0] neuron_0_add, neuron_1_add, neuron_2_add, neuron_3_add, neuron_4_add;
reg [25:0] neuron_5_add, neuron_6_add, neuron_7_add, neuron_8_add, neuron_9_add;
always @(posedge clk) begin
  if(globalreset) begin
    neuron_0_add <= 0;
	neuron_1_add <= 0;
	neuron_2_add <= 0;
	neuron_3_add <= 0;
	neuron_4_add <= 0;
	neuron_5_add <= 0;
	neuron_6_add <= 0;
	neuron_7_add <= 0;
	neuron_8_add <= 0;
	neuron_9_add <= 0;
  end
  else begin
    if(N >= 11) begin  // Maybe 12 or 13, check waveforms for sure
	  neuron_0_add <= neuron_0_add + neuron_0_add_27_out;
	  neuron_1_add <= neuron_1_add + neuron_1_add_27_out;
	  neuron_2_add <= neuron_2_add + neuron_2_add_27_out;
	  neuron_3_add <= neuron_3_add + neuron_3_add_27_out;
	  neuron_4_add <= neuron_4_add + neuron_4_add_27_out;
	  neuron_5_add <= neuron_5_add + neuron_5_add_27_out;
	  neuron_6_add <= neuron_6_add + neuron_6_add_27_out;
	  neuron_7_add <= neuron_7_add + neuron_7_add_27_out;
	  neuron_8_add <= neuron_8_add + neuron_8_add_27_out;
	  neuron_9_add <= neuron_9_add + neuron_9_add_27_out;
	end
	else begin
	  neuron_0_add <= 0;
	  neuron_1_add <= 0;
	  neuron_2_add <= 0;
	  neuron_3_add <= 0;
	  neuron_4_add <= 0;
	  neuron_5_add <= 0;
	  neuron_6_add <= 0;
	  neuron_7_add <= 0;
	  neuron_8_add <= 0;
	  neuron_9_add <= 0;
	end
  end
end

// Mapping neurons' outputs to positive numbers and compare them as unsigned numbers
// Work when neurons' outputs have no overflow
wire [25:0] neuron_0_out, neuron_1_out, neuron_2_out, neuron_3_out, neuron_4_out;
wire [25:0] neuron_5_out, neuron_6_out, neuron_7_out, neuron_8_out, neuron_9_out;
assign neuron_0_out = {~neuron_0_add[25], neuron_0_add[24:0]};
assign neuron_1_out = {~neuron_1_add[25], neuron_1_add[24:0]};
assign neuron_2_out = {~neuron_2_add[25], neuron_2_add[24:0]};
assign neuron_3_out = {~neuron_3_add[25], neuron_3_add[24:0]};
assign neuron_4_out = {~neuron_4_add[25], neuron_4_add[24:0]};
assign neuron_5_out = {~neuron_5_add[25], neuron_5_add[24:0]};
assign neuron_6_out = {~neuron_6_add[25], neuron_6_add[24:0]};
assign neuron_7_out = {~neuron_7_add[25], neuron_7_add[24:0]};
assign neuron_8_out = {~neuron_8_add[25], neuron_8_add[24:0]};
assign neuron_9_out = {~neuron_9_add[25], neuron_9_add[24:0]};

// Compare mapping results and determine Image_Number
// Have to do it in parallel to save time. Already use a lot of circuit area. Acceptable to use some more.
// Sequential version: About 10 clock cycles delay.
reg [3:0] max_out;
reg [25:0] max_neuron_out;
reg [25:0] neuron_out [0:9];
neuron_out[0] = neuron_0_out;
neuron_out[1] = neuron_1_out;
neuron_out[2] = neuron_2_out;
neuron_out[3] = neuron_3_out;
neuron_out[4] = neuron_4_out;
neuron_out[5] = neuron_5_out;
neuron_out[6] = neuron_6_out;
neuron_out[7] = neuron_7_out;
neuron_out[8] = neuron_8_out;
neuron_out[9] = neuron_9_out;
always @(posedge clk) begin  // max_out is the index of the output reg.
  if(globalreset) begin
    max_out <= 0;
	max_neuron_out <= 0;
  end
  else begin
    if (N >= 39 && max_out < 10) begin // Threhold value is to be decided
  	  if (max_neuron_out < neuron_out[max_out]) begin
  	      max_neuron_out <= neuron_out[max_out];
  		    Image_Number <= max_out;
  	  end
  	  else
  	    max_neuron_out <= max_neuron_out;
  	  max_out <= max_out + 1;
    end
  	else begin
  	  max_out <= 0
  	  max_neuron_out <= 0;
  	end
  end
end

always @(posedge clk) begin
  if(globalreset) begin
    Output_Valid <= 0;
  end
  else begin
    if(max_out == 10)  // Output_Valid only asserts only one clock cycle. It should be enough.
	  Output_Valid <= 1;
  	else
  	  Output_Valid <= 0;
  end
end
/*
// Parallel version. Not sure if it can work. About 5 clock cycles delay.
// Image_Number and Output_Valid are wire signals in this case
Max_10 max_10(
.neuron_clk,
.globalreset,
.N,
.neuron_0_out,
.neuron_1_out,
.neuron_2_out,
.neuron_3_out,
.neuron_4_out,
.neuron_5_out,
.neuron_6_out,
.neuron_7_out,
.neuron_8_out,
.neuron_9_out,
.Output_Valid,
.Image_Number
);  */

endmodule
/*
// A main problem for parallel solution is how to determine the location of the largest number.
module Max_10(
input clk,
input GlobalReset,
input N,
input [25:0] Max_in_0,
input [25:0] Max_in_1,
input [25:0] Max_in_2,
input [25:0] Max_in_3,
input [25:0] Max_in_4,
input [25:0] Max_in_5,
input [25:0] Max_in_6,
input [25:0] Max_in_7,
input [25:0] Max_in_8,
input [25:0] Max_in_9,
output reg output_valid,
output reg [3:0] Max_out
);

reg [25:0] comparator_0, comparator_1, comparator_2, comparator_3, comparator_4, comparator_5;
reg [25:0] comparator_6, comparator_7, comparator_8, comparator_9, comparator_10;
always @(posedge clk) begin
  if(GlobalReset)
    Max_out <= 0;
	output_valid <= 0;
	comparator_0 <= 0;
	comparator_1 <= 0;
	comparator_2 <= 0;
	comparator_3 <= 0;
	comparator_4 <= 0;
	comparator_5 <= 0;
	comparator_6 <= 0;
	comparator_7 <= 0;
	comparator_8 <= 0;
	comparator_9 <= 0;
	comparator_10 <= 0;
  else begin
    if(N >= 43 && (!output_valid)) begin
	  case(comparator_10):  // Or use if statement
	    Max_in_0: Max_out <= 0;
		Max_in_1: Max_out <= 1;
		Max_in_2: Max_out <= 2;
		Max_in_3: Max_out <= 3;
		Max_in_4: Max_out <= 4;
		Max_in_5: Max_out <= 5;
		Max_in_6: Max_out <= 6;
		Max_in_7: Max_out <= 7;
		Max_in_8: Max_out <= 8;
		Max_in_9: Max_out <= 9;
		default: Max_out <= 0;
	  endcase
	  output_valid <= 1;
	end
    else if(N >= 39 && (!output_valid)) begin
	  if(Max_in_0 > Max_in_1)
	    comparator_0 <= Max_in_0;
	  else
	    comparator_0 <= Max_in_1;
	  if(Max_in_2 > Max_in_3)
	    comparator_1 <= Max_in_2;
	  else
	    comparator_1 <= Max_in_3;
	  if(Max_in_4 > Max_in_5)
	    comparator_2 <= Max_in_4;
	  else
	    comparator_2 <= Max_in_5;
	  if(Max_in_6 > Max_in_7)
	    comparator_3 <= Max_in_6;
	  else
	    comparator_3 <= Max_in_7;
	  if(Max_in_8 > Max_in_9)
	    comparator_4 <= Max_in_8;
	  else
	    comparator_4 <= Max_in_9;
	  if(comparator_0 > comparator_1)
	    comparator_5 <= comparator_0;
	  else
	    comparator_5 <= comparator_1;
	  if(comparator_2 > comparator_3)
	    comparator_6 <= comparator_2;
	  else
	    comparator_6 <= comparator_3;
	  comparator_7 <= comparator_4;
	  if(comparator_5 > comparator_6)
	    comparator_8 <= comparator_5;
	  else
	    comparator_8 <= comparator_6;
	  comparator_9 <= comparator_7;
	  if(comparator_8 > comparator_9)
	    comparator_10 <= comparator_8;
	  else
	    comparator_10 <= comparator_9;
	end
	else begin
	  Max_out <= 0;
	  output_valid <= 0;
	  comparator_0 <= 0;
	  comparator_1 <= 0;
	  comparator_2 <= 0;
	  comparator_3 <= 0;
	  comparator_4 <= 0;
	  comparator_5 <= 0;
	  comparator_6 <= 0;
	  comparator_7 <= 0;
	  comparator_8 <= 0;
	  comparator_9 <= 0;
	  comparator_10 <= 0;
	end
  end
end

endmodule
